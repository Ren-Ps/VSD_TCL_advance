
module openMSP430(aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dmem_addr_0_, dmem_addr_1_, dmem_addr_2_, dmem_addr_3_, dmem_addr_4_, dmem_addr_5_, dmem_addr_6_, dmem_addr_7_, dmem_addr_8_, dmem_addr_9_, dmem_addr_10_, dmem_addr_11_, dmem_addr_12_, dmem_cen
, dmem_din_0_, dmem_din_1_, dmem_din_2_, dmem_din_3_, dmem_din_4_, dmem_din_5_, dmem_din_6_, dmem_din_7_, dmem_din_8_, dmem_din_9_, dmem_din_10_, dmem_din_11_, dmem_din_12_, dmem_din_13_, dmem_din_14_, dmem_din_15_, dmem_wen_0_, dmem_wen_1_, irq_acc_0_, irq_acc_1_, irq_acc_2_
, irq_acc_3_, irq_acc_4_, irq_acc_5_, irq_acc_6_, irq_acc_7_, irq_acc_8_, irq_acc_9_, irq_acc_10_, irq_acc_11_, irq_acc_12_, irq_acc_13_, lfxt_enable, lfxt_wkup, mclk, dma_dout_0_, dma_dout_1_, dma_dout_2_, dma_dout_3_, dma_dout_4_, dma_dout_5_, dma_dout_6_
, dma_dout_7_, dma_dout_8_, dma_dout_9_, dma_dout_10_, dma_dout_11_, dma_dout_12_, dma_dout_13_, dma_dout_14_, dma_dout_15_, dma_ready, dma_resp, per_addr_0_, per_addr_1_, per_addr_2_, per_addr_3_, per_addr_4_, per_addr_5_, per_addr_6_, per_addr_7_, per_addr_8_, per_addr_9_
, per_addr_10_, per_addr_11_, per_addr_12_, per_addr_13_, per_din_0_, per_din_1_, per_din_2_, per_din_3_, per_din_4_, per_din_5_, per_din_6_, per_din_7_, per_din_8_, per_din_9_, per_din_10_, per_din_11_, per_din_12_, per_din_13_, per_din_14_, per_din_15_, per_en
, per_we_0_, per_we_1_, pmem_addr_0_, pmem_addr_1_, pmem_addr_2_, pmem_addr_3_, pmem_addr_4_, pmem_addr_5_, pmem_addr_6_, pmem_addr_7_, pmem_addr_8_, pmem_addr_9_, pmem_addr_10_, pmem_addr_11_, pmem_addr_12_, pmem_addr_13_, pmem_cen, pmem_din_0_, pmem_din_1_, pmem_din_2_, pmem_din_3_
, pmem_din_4_, pmem_din_5_, pmem_din_6_, pmem_din_7_, pmem_din_8_, pmem_din_9_, pmem_din_10_, pmem_din_11_, pmem_din_12_, pmem_din_13_, pmem_din_14_, pmem_din_15_, pmem_wen_0_, pmem_wen_1_, puc_rst, smclk, smclk_en, cpu_en, dbg_en, dbg_i2c_addr_0_, dbg_i2c_addr_1_
, dbg_i2c_addr_2_, dbg_i2c_addr_3_, dbg_i2c_addr_4_, dbg_i2c_addr_5_, dbg_i2c_addr_6_, dbg_i2c_broadcast_0_, dbg_i2c_broadcast_1_, dbg_i2c_broadcast_2_, dbg_i2c_broadcast_3_, dbg_i2c_broadcast_4_, dbg_i2c_broadcast_5_, dbg_i2c_broadcast_6_, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dmem_dout_0_, dmem_dout_1_, dmem_dout_2_, dmem_dout_3_, dmem_dout_4_
, dmem_dout_5_, dmem_dout_6_, dmem_dout_7_, dmem_dout_8_, dmem_dout_9_, dmem_dout_10_, dmem_dout_11_, dmem_dout_12_, dmem_dout_13_, dmem_dout_14_, dmem_dout_15_, irq_0_, irq_1_, irq_2_, irq_3_, irq_4_, irq_5_, irq_6_, irq_7_, irq_8_, irq_9_
, irq_10_, irq_11_, irq_12_, irq_13_, lfxt_clk, dma_addr_1_, dma_addr_2_, dma_addr_3_, dma_addr_4_, dma_addr_5_, dma_addr_6_, dma_addr_7_, dma_addr_8_, dma_addr_9_, dma_addr_10_, dma_addr_11_, dma_addr_12_, dma_addr_13_, dma_addr_14_, dma_addr_15_, dma_din_0_
, dma_din_1_, dma_din_2_, dma_din_3_, dma_din_4_, dma_din_5_, dma_din_6_, dma_din_7_, dma_din_8_, dma_din_9_, dma_din_10_, dma_din_11_, dma_din_12_, dma_din_13_, dma_din_14_, dma_din_15_, dma_en, dma_priority, dma_we_0_, dma_we_1_, dma_wkup, nmi
, per_dout_0_, per_dout_1_, per_dout_2_, per_dout_3_, per_dout_4_, per_dout_5_, per_dout_6_, per_dout_7_, per_dout_8_, per_dout_9_, per_dout_10_, per_dout_11_, per_dout_12_, per_dout_13_, per_dout_14_, per_dout_15_, pmem_dout_0_, pmem_dout_1_, pmem_dout_2_, pmem_dout_3_, pmem_dout_4_
, pmem_dout_5_, pmem_dout_6_, pmem_dout_7_, pmem_dout_8_, pmem_dout_9_, pmem_dout_10_, pmem_dout_11_, pmem_dout_12_, pmem_dout_13_, pmem_dout_14_, pmem_dout_15_, reset_n, scan_enable, scan_mode, wkup);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  output aclk;
  wire aclk;
  output aclk_en;
  wire aclk_en;
  wire  clock_module_0.UNUSED_cpuoff ;
  wire  clock_module_0.aclk_div_0_ ;
  wire  clock_module_0.aclk_div_1_ ;
  wire  clock_module_0.aclk_div_2_ ;
  wire  clock_module_0.bcsctl1_4_ ;
  wire  clock_module_0.bcsctl1_5_ ;
  wire  clock_module_0.bcsctl1_rd_12_ ;
  wire  clock_module_0.bcsctl1_rd_13_ ;
  wire  clock_module_0.bcsctl2_1_ ;
  wire  clock_module_0.bcsctl2_2_ ;
  wire  clock_module_0.bcsctl2_3_ ;
  wire  clock_module_0.bcsctl2_rd_1_ ;
  wire  clock_module_0.bcsctl2_rd_2_ ;
  wire  clock_module_0.bcsctl2_rd_3_ ;
  wire  clock_module_0.dbg_cpu_reset ;
  wire  clock_module_0.dbg_rst ;
  wire  clock_module_0.dbg_rst_nxt ;
  wire  clock_module_0.lfxt_clk_dly ;
  wire  clock_module_0.lfxt_clk_s ;
  wire  clock_module_0.oscoff ;
  wire  clock_module_0.por ;
  wire  clock_module_0.por_a ;
  wire  clock_module_0.puc_a ;
  wire  clock_module_0.puc_noscan_n ;
  wire  clock_module_0.scg1 ;
  wire  clock_module_0.smclk_div_0_ ;
  wire  clock_module_0.smclk_div_1_ ;
  wire  clock_module_0.smclk_div_2_ ;
  wire  clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ;
  wire  clock_module_0.sync_cell_puc.data_in ;
  wire  clock_module_0.sync_cell_puc.data_sync_0_ ;
  wire  clock_module_0.sync_reset_por.data_sync_0_ ;
  wire  clock_module_0.wdt_reset ;
  input cpu_en;
  wire cpu_en;
  wire  dbg_0.UNUSED_eu_mab_0_ ;
  wire  dbg_0.UNUSED_eu_mab_10_ ;
  wire  dbg_0.UNUSED_eu_mab_11_ ;
  wire  dbg_0.UNUSED_eu_mab_12_ ;
  wire  dbg_0.UNUSED_eu_mab_13_ ;
  wire  dbg_0.UNUSED_eu_mab_14_ ;
  wire  dbg_0.UNUSED_eu_mab_15_ ;
  wire  dbg_0.UNUSED_eu_mab_1_ ;
  wire  dbg_0.UNUSED_eu_mab_2_ ;
  wire  dbg_0.UNUSED_eu_mab_3_ ;
  wire  dbg_0.UNUSED_eu_mab_4_ ;
  wire  dbg_0.UNUSED_eu_mab_5_ ;
  wire  dbg_0.UNUSED_eu_mab_6_ ;
  wire  dbg_0.UNUSED_eu_mab_7_ ;
  wire  dbg_0.UNUSED_eu_mab_8_ ;
  wire  dbg_0.UNUSED_eu_mab_9_ ;
  wire  dbg_0.UNUSED_eu_mb_en ;
  wire  dbg_0.UNUSED_eu_mb_wr_0_ ;
  wire  dbg_0.UNUSED_eu_mb_wr_1_ ;
  wire  dbg_0.UNUSED_pc_0_ ;
  wire  dbg_0.UNUSED_pc_10_ ;
  wire  dbg_0.UNUSED_pc_11_ ;
  wire  dbg_0.UNUSED_pc_12_ ;
  wire  dbg_0.UNUSED_pc_13_ ;
  wire  dbg_0.UNUSED_pc_14_ ;
  wire  dbg_0.UNUSED_pc_15_ ;
  wire  dbg_0.UNUSED_pc_1_ ;
  wire  dbg_0.UNUSED_pc_2_ ;
  wire  dbg_0.UNUSED_pc_3_ ;
  wire  dbg_0.UNUSED_pc_4_ ;
  wire  dbg_0.UNUSED_pc_5_ ;
  wire  dbg_0.UNUSED_pc_6_ ;
  wire  dbg_0.UNUSED_pc_7_ ;
  wire  dbg_0.UNUSED_pc_8_ ;
  wire  dbg_0.UNUSED_pc_9_ ;
  wire  dbg_0.cpu_ctl_3_ ;
  wire  dbg_0.cpu_ctl_4_ ;
  wire  dbg_0.cpu_ctl_5_ ;
  wire  dbg_0.cpu_stat_2_ ;
  wire  dbg_0.cpu_stat_3_ ;
  wire  dbg_0.cpu_stat_full_0_ ;
  wire  dbg_0.dbg_addr_0_ ;
  wire  dbg_0.dbg_addr_1_ ;
  wire  dbg_0.dbg_addr_2_ ;
  wire  dbg_0.dbg_addr_3_ ;
  wire  dbg_0.dbg_addr_4_ ;
  wire  dbg_0.dbg_addr_5_ ;
  wire  dbg_0.dbg_din_0_ ;
  wire  dbg_0.dbg_din_10_ ;
  wire  dbg_0.dbg_din_11_ ;
  wire  dbg_0.dbg_din_12_ ;
  wire  dbg_0.dbg_din_13_ ;
  wire  dbg_0.dbg_din_14_ ;
  wire  dbg_0.dbg_din_15_ ;
  wire  dbg_0.dbg_din_1_ ;
  wire  dbg_0.dbg_din_2_ ;
  wire  dbg_0.dbg_din_3_ ;
  wire  dbg_0.dbg_din_4_ ;
  wire  dbg_0.dbg_din_5_ ;
  wire  dbg_0.dbg_din_6_ ;
  wire  dbg_0.dbg_din_7_ ;
  wire  dbg_0.dbg_din_8_ ;
  wire  dbg_0.dbg_din_9_ ;
  wire  dbg_0.dbg_dout_0_ ;
  wire  dbg_0.dbg_dout_10_ ;
  wire  dbg_0.dbg_dout_11_ ;
  wire  dbg_0.dbg_dout_12_ ;
  wire  dbg_0.dbg_dout_13_ ;
  wire  dbg_0.dbg_dout_14_ ;
  wire  dbg_0.dbg_dout_15_ ;
  wire  dbg_0.dbg_dout_1_ ;
  wire  dbg_0.dbg_dout_2_ ;
  wire  dbg_0.dbg_dout_3_ ;
  wire  dbg_0.dbg_dout_4_ ;
  wire  dbg_0.dbg_dout_5_ ;
  wire  dbg_0.dbg_dout_6_ ;
  wire  dbg_0.dbg_dout_7_ ;
  wire  dbg_0.dbg_dout_8_ ;
  wire  dbg_0.dbg_dout_9_ ;
  wire  dbg_0.dbg_halt_cmd ;
  wire  dbg_0.dbg_i2c_0.dbg_bw ;
  wire  dbg_0.dbg_i2c_0.dbg_rd ;
  wire  dbg_0.dbg_i2c_0.dbg_state_0_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_1_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_2_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_0_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_1_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_2_ ;
  wire  dbg_0.dbg_i2c_0.dbg_wr ;
  wire  dbg_0.dbg_i2c_0.i2c_active_seq ;
  wire  dbg_0.dbg_i2c_0.i2c_state_0_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_1_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_2_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_0_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_1_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ;
  wire  dbg_0.dbg_i2c_0.mem_burst ;
  wire  dbg_0.dbg_i2c_0.mem_burst_end ;
  wire  dbg_0.dbg_i2c_0.mem_burst_rd ;
  wire  dbg_0.dbg_i2c_0.mem_burst_wr ;
  wire  dbg_0.dbg_i2c_0.mem_bw ;
  wire  dbg_0.dbg_i2c_0.scl ;
  wire  dbg_0.dbg_i2c_0.scl_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.scl_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.scl_dly ;
  wire  dbg_0.dbg_i2c_0.scl_re ;
  wire  dbg_0.dbg_i2c_0.scl_re_dly_0_ ;
  wire  dbg_0.dbg_i2c_0.scl_re_dly_1_ ;
  wire  dbg_0.dbg_i2c_0.scl_sync ;
  wire  dbg_0.dbg_i2c_0.scl_sync_n ;
  wire  dbg_0.dbg_i2c_0.sda_in ;
  wire  dbg_0.dbg_i2c_0.sda_in_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.sda_in_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.sda_in_dly ;
  wire  dbg_0.dbg_i2c_0.sda_in_sync ;
  wire  dbg_0.dbg_i2c_0.sda_in_sync_n ;
  wire  dbg_0.dbg_i2c_0.shift_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_2_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_3_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_4_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_5_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_6_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_7_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_8_ ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ;
  wire  dbg_0.dbg_mem_addr_0_ ;
  wire  dbg_0.dbg_mem_addr_10_ ;
  wire  dbg_0.dbg_mem_addr_11_ ;
  wire  dbg_0.dbg_mem_addr_12_ ;
  wire  dbg_0.dbg_mem_addr_13_ ;
  wire  dbg_0.dbg_mem_addr_14_ ;
  wire  dbg_0.dbg_mem_addr_15_ ;
  wire  dbg_0.dbg_mem_addr_1_ ;
  wire  dbg_0.dbg_mem_addr_2_ ;
  wire  dbg_0.dbg_mem_addr_3_ ;
  wire  dbg_0.dbg_mem_addr_4_ ;
  wire  dbg_0.dbg_mem_addr_5_ ;
  wire  dbg_0.dbg_mem_addr_6_ ;
  wire  dbg_0.dbg_mem_addr_7_ ;
  wire  dbg_0.dbg_mem_addr_8_ ;
  wire  dbg_0.dbg_mem_addr_9_ ;
  wire  dbg_0.dbg_mem_din_0_ ;
  wire  dbg_0.dbg_mem_din_10_ ;
  wire  dbg_0.dbg_mem_din_11_ ;
  wire  dbg_0.dbg_mem_din_12_ ;
  wire  dbg_0.dbg_mem_din_13_ ;
  wire  dbg_0.dbg_mem_din_14_ ;
  wire  dbg_0.dbg_mem_din_15_ ;
  wire  dbg_0.dbg_mem_din_1_ ;
  wire  dbg_0.dbg_mem_din_2_ ;
  wire  dbg_0.dbg_mem_din_3_ ;
  wire  dbg_0.dbg_mem_din_4_ ;
  wire  dbg_0.dbg_mem_din_5_ ;
  wire  dbg_0.dbg_mem_din_6_ ;
  wire  dbg_0.dbg_mem_din_7_ ;
  wire  dbg_0.dbg_mem_din_8_ ;
  wire  dbg_0.dbg_mem_din_9_ ;
  wire  dbg_0.dbg_mem_en ;
  wire  dbg_0.dbg_mem_rd ;
  wire  dbg_0.dbg_mem_rd_dly ;
  wire  dbg_0.dbg_mem_wr_0_ ;
  wire  dbg_0.dbg_mem_wr_1_ ;
  wire  dbg_0.dbg_rd_rdy ;
  wire  dbg_0.dbg_reg_din_0_ ;
  wire  dbg_0.dbg_reg_din_10_ ;
  wire  dbg_0.dbg_reg_din_11_ ;
  wire  dbg_0.dbg_reg_din_12_ ;
  wire  dbg_0.dbg_reg_din_13_ ;
  wire  dbg_0.dbg_reg_din_14_ ;
  wire  dbg_0.dbg_reg_din_15_ ;
  wire  dbg_0.dbg_reg_din_1_ ;
  wire  dbg_0.dbg_reg_din_2_ ;
  wire  dbg_0.dbg_reg_din_3_ ;
  wire  dbg_0.dbg_reg_din_4_ ;
  wire  dbg_0.dbg_reg_din_5_ ;
  wire  dbg_0.dbg_reg_din_6_ ;
  wire  dbg_0.dbg_reg_din_7_ ;
  wire  dbg_0.dbg_reg_din_8_ ;
  wire  dbg_0.dbg_reg_din_9_ ;
  wire  dbg_0.dbg_reg_wr ;
  wire  dbg_0.decode_noirq ;
  wire  dbg_0.fe_mdb_in_0_ ;
  wire  dbg_0.fe_mdb_in_10_ ;
  wire  dbg_0.fe_mdb_in_11_ ;
  wire  dbg_0.fe_mdb_in_12_ ;
  wire  dbg_0.fe_mdb_in_13_ ;
  wire  dbg_0.fe_mdb_in_14_ ;
  wire  dbg_0.fe_mdb_in_15_ ;
  wire  dbg_0.fe_mdb_in_1_ ;
  wire  dbg_0.fe_mdb_in_2_ ;
  wire  dbg_0.fe_mdb_in_3_ ;
  wire  dbg_0.fe_mdb_in_4_ ;
  wire  dbg_0.fe_mdb_in_5_ ;
  wire  dbg_0.fe_mdb_in_6_ ;
  wire  dbg_0.fe_mdb_in_7_ ;
  wire  dbg_0.fe_mdb_in_8_ ;
  wire  dbg_0.fe_mdb_in_9_ ;
  wire  dbg_0.halt_flag ;
  wire  dbg_0.inc_step_0_ ;
  wire  dbg_0.inc_step_1_ ;
  wire  dbg_0.istep ;
  wire  dbg_0.mem_cnt_0_ ;
  wire  dbg_0.mem_cnt_10_ ;
  wire  dbg_0.mem_cnt_11_ ;
  wire  dbg_0.mem_cnt_12_ ;
  wire  dbg_0.mem_cnt_13_ ;
  wire  dbg_0.mem_cnt_14_ ;
  wire  dbg_0.mem_cnt_15_ ;
  wire  dbg_0.mem_cnt_1_ ;
  wire  dbg_0.mem_cnt_2_ ;
  wire  dbg_0.mem_cnt_3_ ;
  wire  dbg_0.mem_cnt_4_ ;
  wire  dbg_0.mem_cnt_5_ ;
  wire  dbg_0.mem_cnt_6_ ;
  wire  dbg_0.mem_cnt_7_ ;
  wire  dbg_0.mem_cnt_8_ ;
  wire  dbg_0.mem_cnt_9_ ;
  wire  dbg_0.mem_ctl_1_ ;
  wire  dbg_0.mem_ctl_2_ ;
  wire  dbg_0.mem_data_0_ ;
  wire  dbg_0.mem_data_10_ ;
  wire  dbg_0.mem_data_11_ ;
  wire  dbg_0.mem_data_12_ ;
  wire  dbg_0.mem_data_13_ ;
  wire  dbg_0.mem_data_14_ ;
  wire  dbg_0.mem_data_15_ ;
  wire  dbg_0.mem_data_1_ ;
  wire  dbg_0.mem_data_2_ ;
  wire  dbg_0.mem_data_3_ ;
  wire  dbg_0.mem_data_4_ ;
  wire  dbg_0.mem_data_5_ ;
  wire  dbg_0.mem_data_6_ ;
  wire  dbg_0.mem_data_7_ ;
  wire  dbg_0.mem_data_8_ ;
  wire  dbg_0.mem_data_9_ ;
  wire  dbg_0.mem_start ;
  wire  dbg_0.mem_startb ;
  wire  dbg_0.mem_state_0_ ;
  wire  dbg_0.mem_state_1_ ;
  wire  dbg_0.mem_state_nxt_0_ ;
  wire  dbg_0.mem_state_nxt_1_ ;
  input dbg_en;
  wire dbg_en;
  output dbg_freeze;
  wire dbg_freeze;
  input dbg_i2c_addr_0_;
  wire dbg_i2c_addr_0_;
  input dbg_i2c_addr_1_;
  wire dbg_i2c_addr_1_;
  input dbg_i2c_addr_2_;
  wire dbg_i2c_addr_2_;
  input dbg_i2c_addr_3_;
  wire dbg_i2c_addr_3_;
  input dbg_i2c_addr_4_;
  wire dbg_i2c_addr_4_;
  input dbg_i2c_addr_5_;
  wire dbg_i2c_addr_5_;
  input dbg_i2c_addr_6_;
  wire dbg_i2c_addr_6_;
  input dbg_i2c_broadcast_0_;
  wire dbg_i2c_broadcast_0_;
  input dbg_i2c_broadcast_1_;
  wire dbg_i2c_broadcast_1_;
  input dbg_i2c_broadcast_2_;
  wire dbg_i2c_broadcast_2_;
  input dbg_i2c_broadcast_3_;
  wire dbg_i2c_broadcast_3_;
  input dbg_i2c_broadcast_4_;
  wire dbg_i2c_broadcast_4_;
  input dbg_i2c_broadcast_5_;
  wire dbg_i2c_broadcast_5_;
  input dbg_i2c_broadcast_6_;
  wire dbg_i2c_broadcast_6_;
  input dbg_i2c_scl;
  wire dbg_i2c_scl;
  input dbg_i2c_sda_in;
  wire dbg_i2c_sda_in;
  output dbg_i2c_sda_out;
  wire dbg_i2c_sda_out;
  input dbg_uart_rxd;
  wire dbg_uart_rxd;
  output dbg_uart_txd;
  wire dbg_uart_txd;
  input dco_clk;
  wire dco_clk;
  output dco_enable;
  wire dco_enable;
  output dco_wkup;
  wire dco_wkup;
  input dma_addr_10_;
  wire dma_addr_10_;
  input dma_addr_11_;
  wire dma_addr_11_;
  input dma_addr_12_;
  wire dma_addr_12_;
  input dma_addr_13_;
  wire dma_addr_13_;
  input dma_addr_14_;
  wire dma_addr_14_;
  input dma_addr_15_;
  wire dma_addr_15_;
  input dma_addr_1_;
  wire dma_addr_1_;
  input dma_addr_2_;
  wire dma_addr_2_;
  input dma_addr_3_;
  wire dma_addr_3_;
  input dma_addr_4_;
  wire dma_addr_4_;
  input dma_addr_5_;
  wire dma_addr_5_;
  input dma_addr_6_;
  wire dma_addr_6_;
  input dma_addr_7_;
  wire dma_addr_7_;
  input dma_addr_8_;
  wire dma_addr_8_;
  input dma_addr_9_;
  wire dma_addr_9_;
  input dma_din_0_;
  wire dma_din_0_;
  input dma_din_10_;
  wire dma_din_10_;
  input dma_din_11_;
  wire dma_din_11_;
  input dma_din_12_;
  wire dma_din_12_;
  input dma_din_13_;
  wire dma_din_13_;
  input dma_din_14_;
  wire dma_din_14_;
  input dma_din_15_;
  wire dma_din_15_;
  input dma_din_1_;
  wire dma_din_1_;
  input dma_din_2_;
  wire dma_din_2_;
  input dma_din_3_;
  wire dma_din_3_;
  input dma_din_4_;
  wire dma_din_4_;
  input dma_din_5_;
  wire dma_din_5_;
  input dma_din_6_;
  wire dma_din_6_;
  input dma_din_7_;
  wire dma_din_7_;
  input dma_din_8_;
  wire dma_din_8_;
  input dma_din_9_;
  wire dma_din_9_;
  output dma_dout_0_;
  wire dma_dout_0_;
  output dma_dout_10_;
  wire dma_dout_10_;
  output dma_dout_11_;
  wire dma_dout_11_;
  output dma_dout_12_;
  wire dma_dout_12_;
  output dma_dout_13_;
  wire dma_dout_13_;
  output dma_dout_14_;
  wire dma_dout_14_;
  output dma_dout_15_;
  wire dma_dout_15_;
  output dma_dout_1_;
  wire dma_dout_1_;
  output dma_dout_2_;
  wire dma_dout_2_;
  output dma_dout_3_;
  wire dma_dout_3_;
  output dma_dout_4_;
  wire dma_dout_4_;
  output dma_dout_5_;
  wire dma_dout_5_;
  output dma_dout_6_;
  wire dma_dout_6_;
  output dma_dout_7_;
  wire dma_dout_7_;
  output dma_dout_8_;
  wire dma_dout_8_;
  output dma_dout_9_;
  wire dma_dout_9_;
  input dma_en;
  wire dma_en;
  input dma_priority;
  wire dma_priority;
  output dma_ready;
  wire dma_ready;
  output dma_resp;
  wire dma_resp;
  input dma_we_0_;
  wire dma_we_0_;
  input dma_we_1_;
  wire dma_we_1_;
  input dma_wkup;
  wire dma_wkup;
  output dmem_addr_0_;
  wire dmem_addr_0_;
  output dmem_addr_10_;
  wire dmem_addr_10_;
  output dmem_addr_11_;
  wire dmem_addr_11_;
  output dmem_addr_12_;
  wire dmem_addr_12_;
  output dmem_addr_1_;
  wire dmem_addr_1_;
  output dmem_addr_2_;
  wire dmem_addr_2_;
  output dmem_addr_3_;
  wire dmem_addr_3_;
  output dmem_addr_4_;
  wire dmem_addr_4_;
  output dmem_addr_5_;
  wire dmem_addr_5_;
  output dmem_addr_6_;
  wire dmem_addr_6_;
  output dmem_addr_7_;
  wire dmem_addr_7_;
  output dmem_addr_8_;
  wire dmem_addr_8_;
  output dmem_addr_9_;
  wire dmem_addr_9_;
  output dmem_cen;
  wire dmem_cen;
  output dmem_din_0_;
  wire dmem_din_0_;
  output dmem_din_10_;
  wire dmem_din_10_;
  output dmem_din_11_;
  wire dmem_din_11_;
  output dmem_din_12_;
  wire dmem_din_12_;
  output dmem_din_13_;
  wire dmem_din_13_;
  output dmem_din_14_;
  wire dmem_din_14_;
  output dmem_din_15_;
  wire dmem_din_15_;
  output dmem_din_1_;
  wire dmem_din_1_;
  output dmem_din_2_;
  wire dmem_din_2_;
  output dmem_din_3_;
  wire dmem_din_3_;
  output dmem_din_4_;
  wire dmem_din_4_;
  output dmem_din_5_;
  wire dmem_din_5_;
  output dmem_din_6_;
  wire dmem_din_6_;
  output dmem_din_7_;
  wire dmem_din_7_;
  output dmem_din_8_;
  wire dmem_din_8_;
  output dmem_din_9_;
  wire dmem_din_9_;
  input dmem_dout_0_;
  wire dmem_dout_0_;
  input dmem_dout_10_;
  wire dmem_dout_10_;
  input dmem_dout_11_;
  wire dmem_dout_11_;
  input dmem_dout_12_;
  wire dmem_dout_12_;
  input dmem_dout_13_;
  wire dmem_dout_13_;
  input dmem_dout_14_;
  wire dmem_dout_14_;
  input dmem_dout_15_;
  wire dmem_dout_15_;
  input dmem_dout_1_;
  wire dmem_dout_1_;
  input dmem_dout_2_;
  wire dmem_dout_2_;
  input dmem_dout_3_;
  wire dmem_dout_3_;
  input dmem_dout_4_;
  wire dmem_dout_4_;
  input dmem_dout_5_;
  wire dmem_dout_5_;
  input dmem_dout_6_;
  wire dmem_dout_6_;
  input dmem_dout_7_;
  wire dmem_dout_7_;
  input dmem_dout_8_;
  wire dmem_dout_8_;
  input dmem_dout_9_;
  wire dmem_dout_9_;
  output dmem_wen_0_;
  wire dmem_wen_0_;
  output dmem_wen_1_;
  wire dmem_wen_1_;
  wire  execution_unit_0.UNUSED_inst_ad_idx ;
  wire  execution_unit_0.UNUSED_inst_ad_symb ;
  wire  execution_unit_0.alu_0.N ;
  wire  execution_unit_0.alu_0.UNUSED_inst_alu ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_call ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_push ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_reti ;
  wire  execution_unit_0.alu_0.Z ;
  wire  execution_unit_0.alu_0.alu_out_0_ ;
  wire  execution_unit_0.alu_0.alu_out_10_ ;
  wire  execution_unit_0.alu_0.alu_out_11_ ;
  wire  execution_unit_0.alu_0.alu_out_12_ ;
  wire  execution_unit_0.alu_0.alu_out_13_ ;
  wire  execution_unit_0.alu_0.alu_out_14_ ;
  wire  execution_unit_0.alu_0.alu_out_15_ ;
  wire  execution_unit_0.alu_0.alu_out_1_ ;
  wire  execution_unit_0.alu_0.alu_out_2_ ;
  wire  execution_unit_0.alu_0.alu_out_3_ ;
  wire  execution_unit_0.alu_0.alu_out_4_ ;
  wire  execution_unit_0.alu_0.alu_out_5_ ;
  wire  execution_unit_0.alu_0.alu_out_6_ ;
  wire  execution_unit_0.alu_0.alu_out_7_ ;
  wire  execution_unit_0.alu_0.alu_out_8_ ;
  wire  execution_unit_0.alu_0.alu_out_9_ ;
  wire  execution_unit_0.alu_0.alu_shift_0_ ;
  wire  execution_unit_0.alu_0.alu_shift_10_ ;
  wire  execution_unit_0.alu_0.alu_shift_11_ ;
  wire  execution_unit_0.alu_0.alu_shift_12_ ;
  wire  execution_unit_0.alu_0.alu_shift_13_ ;
  wire  execution_unit_0.alu_0.alu_shift_14_ ;
  wire  execution_unit_0.alu_0.alu_shift_1_ ;
  wire  execution_unit_0.alu_0.alu_shift_2_ ;
  wire  execution_unit_0.alu_0.alu_shift_3_ ;
  wire  execution_unit_0.alu_0.alu_shift_4_ ;
  wire  execution_unit_0.alu_0.alu_shift_5_ ;
  wire  execution_unit_0.alu_0.alu_shift_6_ ;
  wire  execution_unit_0.alu_0.alu_shift_8_ ;
  wire  execution_unit_0.alu_0.alu_shift_9_ ;
  wire  execution_unit_0.alu_0.alu_stat_0_ ;
  wire  execution_unit_0.alu_0.alu_stat_3_ ;
  wire  execution_unit_0.alu_0.alu_stat_wr_0_ ;
  wire  execution_unit_0.alu_0.alu_swpb_0_ ;
  wire  execution_unit_0.alu_0.alu_swpb_8_ ;
  wire  execution_unit_0.alu_0.exec_cycle ;
  wire  execution_unit_0.alu_0.inst_alu_0_ ;
  wire  execution_unit_0.alu_0.inst_alu_10_ ;
  wire  execution_unit_0.alu_0.inst_alu_1_ ;
  wire  execution_unit_0.alu_0.inst_alu_2_ ;
  wire  execution_unit_0.alu_0.inst_alu_3_ ;
  wire  execution_unit_0.alu_0.inst_alu_4_ ;
  wire  execution_unit_0.alu_0.inst_alu_5_ ;
  wire  execution_unit_0.alu_0.inst_alu_6_ ;
  wire  execution_unit_0.alu_0.inst_alu_7_ ;
  wire  execution_unit_0.alu_0.inst_alu_8_ ;
  wire  execution_unit_0.alu_0.inst_alu_9_ ;
  wire  execution_unit_0.alu_0.inst_bw ;
  wire  execution_unit_0.alu_0.inst_jmp_0_ ;
  wire  execution_unit_0.alu_0.inst_jmp_1_ ;
  wire  execution_unit_0.alu_0.inst_jmp_2_ ;
  wire  execution_unit_0.alu_0.inst_jmp_3_ ;
  wire  execution_unit_0.alu_0.inst_jmp_4_ ;
  wire  execution_unit_0.alu_0.inst_jmp_5_ ;
  wire  execution_unit_0.alu_0.inst_jmp_6_ ;
  wire  execution_unit_0.alu_0.inst_so_0_ ;
  wire  execution_unit_0.alu_0.inst_so_1_ ;
  wire  execution_unit_0.alu_0.inst_so_3_ ;
  wire  execution_unit_0.alu_0.inst_so_7_ ;
  wire  execution_unit_0.alu_0.op_dst_0_ ;
  wire  execution_unit_0.alu_0.op_dst_10_ ;
  wire  execution_unit_0.alu_0.op_dst_11_ ;
  wire  execution_unit_0.alu_0.op_dst_12_ ;
  wire  execution_unit_0.alu_0.op_dst_13_ ;
  wire  execution_unit_0.alu_0.op_dst_14_ ;
  wire  execution_unit_0.alu_0.op_dst_15_ ;
  wire  execution_unit_0.alu_0.op_dst_1_ ;
  wire  execution_unit_0.alu_0.op_dst_2_ ;
  wire  execution_unit_0.alu_0.op_dst_3_ ;
  wire  execution_unit_0.alu_0.op_dst_4_ ;
  wire  execution_unit_0.alu_0.op_dst_5_ ;
  wire  execution_unit_0.alu_0.op_dst_6_ ;
  wire  execution_unit_0.alu_0.op_dst_7_ ;
  wire  execution_unit_0.alu_0.op_dst_8_ ;
  wire  execution_unit_0.alu_0.op_dst_9_ ;
  wire  execution_unit_0.alu_0.status_0_ ;
  wire  execution_unit_0.alu_0.status_1_ ;
  wire  execution_unit_0.alu_0.status_2_ ;
  wire  execution_unit_0.alu_0.status_3_ ;
  wire  execution_unit_0.e_state_0_ ;
  wire  execution_unit_0.e_state_1_ ;
  wire  execution_unit_0.e_state_2_ ;
  wire  execution_unit_0.e_state_3_ ;
  wire  execution_unit_0.exec_done ;
  wire  execution_unit_0.gie ;
  wire  execution_unit_0.inst_ad_0_ ;
  wire  execution_unit_0.inst_ad_6_ ;
  wire  execution_unit_0.inst_as_0_ ;
  wire  execution_unit_0.inst_as_1_ ;
  wire  execution_unit_0.inst_as_2_ ;
  wire  execution_unit_0.inst_as_3_ ;
  wire  execution_unit_0.inst_as_4_ ;
  wire  execution_unit_0.inst_as_5_ ;
  wire  execution_unit_0.inst_as_6_ ;
  wire  execution_unit_0.inst_as_7_ ;
  wire  execution_unit_0.inst_dest_0_ ;
  wire  execution_unit_0.inst_dest_10_ ;
  wire  execution_unit_0.inst_dest_11_ ;
  wire  execution_unit_0.inst_dest_12_ ;
  wire  execution_unit_0.inst_dest_13_ ;
  wire  execution_unit_0.inst_dest_14_ ;
  wire  execution_unit_0.inst_dest_15_ ;
  wire  execution_unit_0.inst_dest_1_ ;
  wire  execution_unit_0.inst_dest_2_ ;
  wire  execution_unit_0.inst_dest_3_ ;
  wire  execution_unit_0.inst_dest_4_ ;
  wire  execution_unit_0.inst_dest_5_ ;
  wire  execution_unit_0.inst_dest_6_ ;
  wire  execution_unit_0.inst_dest_7_ ;
  wire  execution_unit_0.inst_dest_8_ ;
  wire  execution_unit_0.inst_dest_9_ ;
  wire  execution_unit_0.inst_dext_0_ ;
  wire  execution_unit_0.inst_dext_10_ ;
  wire  execution_unit_0.inst_dext_11_ ;
  wire  execution_unit_0.inst_dext_12_ ;
  wire  execution_unit_0.inst_dext_13_ ;
  wire  execution_unit_0.inst_dext_14_ ;
  wire  execution_unit_0.inst_dext_15_ ;
  wire  execution_unit_0.inst_dext_1_ ;
  wire  execution_unit_0.inst_dext_2_ ;
  wire  execution_unit_0.inst_dext_3_ ;
  wire  execution_unit_0.inst_dext_4_ ;
  wire  execution_unit_0.inst_dext_5_ ;
  wire  execution_unit_0.inst_dext_6_ ;
  wire  execution_unit_0.inst_dext_7_ ;
  wire  execution_unit_0.inst_dext_8_ ;
  wire  execution_unit_0.inst_dext_9_ ;
  wire  execution_unit_0.inst_irq_rst ;
  wire  execution_unit_0.inst_mov ;
  wire  execution_unit_0.inst_sext_0_ ;
  wire  execution_unit_0.inst_sext_10_ ;
  wire  execution_unit_0.inst_sext_11_ ;
  wire  execution_unit_0.inst_sext_12_ ;
  wire  execution_unit_0.inst_sext_13_ ;
  wire  execution_unit_0.inst_sext_14_ ;
  wire  execution_unit_0.inst_sext_15_ ;
  wire  execution_unit_0.inst_sext_1_ ;
  wire  execution_unit_0.inst_sext_2_ ;
  wire  execution_unit_0.inst_sext_3_ ;
  wire  execution_unit_0.inst_sext_4_ ;
  wire  execution_unit_0.inst_sext_5_ ;
  wire  execution_unit_0.inst_sext_6_ ;
  wire  execution_unit_0.inst_sext_7_ ;
  wire  execution_unit_0.inst_sext_8_ ;
  wire  execution_unit_0.inst_sext_9_ ;
  wire  execution_unit_0.inst_src_0_ ;
  wire  execution_unit_0.inst_src_10_ ;
  wire  execution_unit_0.inst_src_11_ ;
  wire  execution_unit_0.inst_src_12_ ;
  wire  execution_unit_0.inst_src_13_ ;
  wire  execution_unit_0.inst_src_14_ ;
  wire  execution_unit_0.inst_src_15_ ;
  wire  execution_unit_0.inst_src_1_ ;
  wire  execution_unit_0.inst_src_2_ ;
  wire  execution_unit_0.inst_src_3_ ;
  wire  execution_unit_0.inst_src_4_ ;
  wire  execution_unit_0.inst_src_5_ ;
  wire  execution_unit_0.inst_src_6_ ;
  wire  execution_unit_0.inst_src_7_ ;
  wire  execution_unit_0.inst_src_8_ ;
  wire  execution_unit_0.inst_src_9_ ;
  wire  execution_unit_0.inst_type_0_ ;
  wire  execution_unit_0.inst_type_1_ ;
  wire  execution_unit_0.inst_type_2_ ;
  wire  execution_unit_0.mab_lsb ;
  wire  execution_unit_0.mdb_in_0_ ;
  wire  execution_unit_0.mdb_in_10_ ;
  wire  execution_unit_0.mdb_in_11_ ;
  wire  execution_unit_0.mdb_in_12_ ;
  wire  execution_unit_0.mdb_in_13_ ;
  wire  execution_unit_0.mdb_in_14_ ;
  wire  execution_unit_0.mdb_in_15_ ;
  wire  execution_unit_0.mdb_in_1_ ;
  wire  execution_unit_0.mdb_in_2_ ;
  wire  execution_unit_0.mdb_in_3_ ;
  wire  execution_unit_0.mdb_in_4_ ;
  wire  execution_unit_0.mdb_in_5_ ;
  wire  execution_unit_0.mdb_in_6_ ;
  wire  execution_unit_0.mdb_in_7_ ;
  wire  execution_unit_0.mdb_in_8_ ;
  wire  execution_unit_0.mdb_in_9_ ;
  wire  execution_unit_0.mdb_in_buf_0_ ;
  wire  execution_unit_0.mdb_in_buf_10_ ;
  wire  execution_unit_0.mdb_in_buf_11_ ;
  wire  execution_unit_0.mdb_in_buf_12_ ;
  wire  execution_unit_0.mdb_in_buf_13_ ;
  wire  execution_unit_0.mdb_in_buf_14_ ;
  wire  execution_unit_0.mdb_in_buf_15_ ;
  wire  execution_unit_0.mdb_in_buf_1_ ;
  wire  execution_unit_0.mdb_in_buf_2_ ;
  wire  execution_unit_0.mdb_in_buf_3_ ;
  wire  execution_unit_0.mdb_in_buf_4_ ;
  wire  execution_unit_0.mdb_in_buf_5_ ;
  wire  execution_unit_0.mdb_in_buf_6_ ;
  wire  execution_unit_0.mdb_in_buf_7_ ;
  wire  execution_unit_0.mdb_in_buf_8_ ;
  wire  execution_unit_0.mdb_in_buf_9_ ;
  wire  execution_unit_0.mdb_in_buf_en ;
  wire  execution_unit_0.mdb_in_buf_valid ;
  wire  execution_unit_0.mdb_out_0_ ;
  wire  execution_unit_0.mdb_out_10_ ;
  wire  execution_unit_0.mdb_out_11_ ;
  wire  execution_unit_0.mdb_out_12_ ;
  wire  execution_unit_0.mdb_out_13_ ;
  wire  execution_unit_0.mdb_out_14_ ;
  wire  execution_unit_0.mdb_out_15_ ;
  wire  execution_unit_0.mdb_out_1_ ;
  wire  execution_unit_0.mdb_out_2_ ;
  wire  execution_unit_0.mdb_out_3_ ;
  wire  execution_unit_0.mdb_out_4_ ;
  wire  execution_unit_0.mdb_out_5_ ;
  wire  execution_unit_0.mdb_out_6_ ;
  wire  execution_unit_0.mdb_out_7_ ;
  wire  execution_unit_0.mdb_out_8_ ;
  wire  execution_unit_0.mdb_out_9_ ;
  wire  execution_unit_0.mdb_out_nxt_10_ ;
  wire  execution_unit_0.mdb_out_nxt_11_ ;
  wire  execution_unit_0.mdb_out_nxt_12_ ;
  wire  execution_unit_0.mdb_out_nxt_13_ ;
  wire  execution_unit_0.mdb_out_nxt_14_ ;
  wire  execution_unit_0.mdb_out_nxt_15_ ;
  wire  execution_unit_0.mdb_out_nxt_8_ ;
  wire  execution_unit_0.mdb_out_nxt_9_ ;
  wire  execution_unit_0.pc_nxt_0_ ;
  wire  execution_unit_0.pc_nxt_10_ ;
  wire  execution_unit_0.pc_nxt_11_ ;
  wire  execution_unit_0.pc_nxt_12_ ;
  wire  execution_unit_0.pc_nxt_13_ ;
  wire  execution_unit_0.pc_nxt_14_ ;
  wire  execution_unit_0.pc_nxt_15_ ;
  wire  execution_unit_0.pc_nxt_1_ ;
  wire  execution_unit_0.pc_nxt_2_ ;
  wire  execution_unit_0.pc_nxt_3_ ;
  wire  execution_unit_0.pc_nxt_4_ ;
  wire  execution_unit_0.pc_nxt_5_ ;
  wire  execution_unit_0.pc_nxt_6_ ;
  wire  execution_unit_0.pc_nxt_7_ ;
  wire  execution_unit_0.pc_nxt_8_ ;
  wire  execution_unit_0.pc_nxt_9_ ;
  wire  execution_unit_0.pc_sw_10_ ;
  wire  execution_unit_0.pc_sw_11_ ;
  wire  execution_unit_0.pc_sw_12_ ;
  wire  execution_unit_0.pc_sw_13_ ;
  wire  execution_unit_0.pc_sw_14_ ;
  wire  execution_unit_0.pc_sw_15_ ;
  wire  execution_unit_0.pc_sw_8_ ;
  wire  execution_unit_0.pc_sw_9_ ;
  wire  execution_unit_0.pc_sw_wr ;
  wire  execution_unit_0.reg_dest_wr ;
  wire  execution_unit_0.reg_incr ;
  wire  execution_unit_0.reg_pc_call ;
  wire  execution_unit_0.reg_sp_wr ;
  wire  execution_unit_0.reg_sr_clr ;
  wire  execution_unit_0.reg_sr_wr ;
  wire  execution_unit_0.reg_src_0_ ;
  wire  execution_unit_0.reg_src_10_ ;
  wire  execution_unit_0.reg_src_11_ ;
  wire  execution_unit_0.reg_src_12_ ;
  wire  execution_unit_0.reg_src_13_ ;
  wire  execution_unit_0.reg_src_14_ ;
  wire  execution_unit_0.reg_src_15_ ;
  wire  execution_unit_0.reg_src_1_ ;
  wire  execution_unit_0.reg_src_2_ ;
  wire  execution_unit_0.reg_src_3_ ;
  wire  execution_unit_0.reg_src_4_ ;
  wire  execution_unit_0.reg_src_5_ ;
  wire  execution_unit_0.reg_src_6_ ;
  wire  execution_unit_0.reg_src_7_ ;
  wire  execution_unit_0.reg_src_8_ ;
  wire  execution_unit_0.reg_src_9_ ;
  wire  execution_unit_0.register_file_0.r10_0_ ;
  wire  execution_unit_0.register_file_0.r10_10_ ;
  wire  execution_unit_0.register_file_0.r10_11_ ;
  wire  execution_unit_0.register_file_0.r10_12_ ;
  wire  execution_unit_0.register_file_0.r10_13_ ;
  wire  execution_unit_0.register_file_0.r10_14_ ;
  wire  execution_unit_0.register_file_0.r10_15_ ;
  wire  execution_unit_0.register_file_0.r10_1_ ;
  wire  execution_unit_0.register_file_0.r10_2_ ;
  wire  execution_unit_0.register_file_0.r10_3_ ;
  wire  execution_unit_0.register_file_0.r10_4_ ;
  wire  execution_unit_0.register_file_0.r10_5_ ;
  wire  execution_unit_0.register_file_0.r10_6_ ;
  wire  execution_unit_0.register_file_0.r10_7_ ;
  wire  execution_unit_0.register_file_0.r10_8_ ;
  wire  execution_unit_0.register_file_0.r10_9_ ;
  wire  execution_unit_0.register_file_0.r11_0_ ;
  wire  execution_unit_0.register_file_0.r11_10_ ;
  wire  execution_unit_0.register_file_0.r11_11_ ;
  wire  execution_unit_0.register_file_0.r11_12_ ;
  wire  execution_unit_0.register_file_0.r11_13_ ;
  wire  execution_unit_0.register_file_0.r11_14_ ;
  wire  execution_unit_0.register_file_0.r11_15_ ;
  wire  execution_unit_0.register_file_0.r11_1_ ;
  wire  execution_unit_0.register_file_0.r11_2_ ;
  wire  execution_unit_0.register_file_0.r11_3_ ;
  wire  execution_unit_0.register_file_0.r11_4_ ;
  wire  execution_unit_0.register_file_0.r11_5_ ;
  wire  execution_unit_0.register_file_0.r11_6_ ;
  wire  execution_unit_0.register_file_0.r11_7_ ;
  wire  execution_unit_0.register_file_0.r11_8_ ;
  wire  execution_unit_0.register_file_0.r11_9_ ;
  wire  execution_unit_0.register_file_0.r12_0_ ;
  wire  execution_unit_0.register_file_0.r12_10_ ;
  wire  execution_unit_0.register_file_0.r12_11_ ;
  wire  execution_unit_0.register_file_0.r12_12_ ;
  wire  execution_unit_0.register_file_0.r12_13_ ;
  wire  execution_unit_0.register_file_0.r12_14_ ;
  wire  execution_unit_0.register_file_0.r12_15_ ;
  wire  execution_unit_0.register_file_0.r12_1_ ;
  wire  execution_unit_0.register_file_0.r12_2_ ;
  wire  execution_unit_0.register_file_0.r12_3_ ;
  wire  execution_unit_0.register_file_0.r12_4_ ;
  wire  execution_unit_0.register_file_0.r12_5_ ;
  wire  execution_unit_0.register_file_0.r12_6_ ;
  wire  execution_unit_0.register_file_0.r12_7_ ;
  wire  execution_unit_0.register_file_0.r12_8_ ;
  wire  execution_unit_0.register_file_0.r12_9_ ;
  wire  execution_unit_0.register_file_0.r13_0_ ;
  wire  execution_unit_0.register_file_0.r13_10_ ;
  wire  execution_unit_0.register_file_0.r13_11_ ;
  wire  execution_unit_0.register_file_0.r13_12_ ;
  wire  execution_unit_0.register_file_0.r13_13_ ;
  wire  execution_unit_0.register_file_0.r13_14_ ;
  wire  execution_unit_0.register_file_0.r13_15_ ;
  wire  execution_unit_0.register_file_0.r13_1_ ;
  wire  execution_unit_0.register_file_0.r13_2_ ;
  wire  execution_unit_0.register_file_0.r13_3_ ;
  wire  execution_unit_0.register_file_0.r13_4_ ;
  wire  execution_unit_0.register_file_0.r13_5_ ;
  wire  execution_unit_0.register_file_0.r13_6_ ;
  wire  execution_unit_0.register_file_0.r13_7_ ;
  wire  execution_unit_0.register_file_0.r13_8_ ;
  wire  execution_unit_0.register_file_0.r13_9_ ;
  wire  execution_unit_0.register_file_0.r14_0_ ;
  wire  execution_unit_0.register_file_0.r14_10_ ;
  wire  execution_unit_0.register_file_0.r14_11_ ;
  wire  execution_unit_0.register_file_0.r14_12_ ;
  wire  execution_unit_0.register_file_0.r14_13_ ;
  wire  execution_unit_0.register_file_0.r14_14_ ;
  wire  execution_unit_0.register_file_0.r14_15_ ;
  wire  execution_unit_0.register_file_0.r14_1_ ;
  wire  execution_unit_0.register_file_0.r14_2_ ;
  wire  execution_unit_0.register_file_0.r14_3_ ;
  wire  execution_unit_0.register_file_0.r14_4_ ;
  wire  execution_unit_0.register_file_0.r14_5_ ;
  wire  execution_unit_0.register_file_0.r14_6_ ;
  wire  execution_unit_0.register_file_0.r14_7_ ;
  wire  execution_unit_0.register_file_0.r14_8_ ;
  wire  execution_unit_0.register_file_0.r14_9_ ;
  wire  execution_unit_0.register_file_0.r15_0_ ;
  wire  execution_unit_0.register_file_0.r15_10_ ;
  wire  execution_unit_0.register_file_0.r15_11_ ;
  wire  execution_unit_0.register_file_0.r15_12_ ;
  wire  execution_unit_0.register_file_0.r15_13_ ;
  wire  execution_unit_0.register_file_0.r15_14_ ;
  wire  execution_unit_0.register_file_0.r15_15_ ;
  wire  execution_unit_0.register_file_0.r15_1_ ;
  wire  execution_unit_0.register_file_0.r15_2_ ;
  wire  execution_unit_0.register_file_0.r15_3_ ;
  wire  execution_unit_0.register_file_0.r15_4_ ;
  wire  execution_unit_0.register_file_0.r15_5_ ;
  wire  execution_unit_0.register_file_0.r15_6_ ;
  wire  execution_unit_0.register_file_0.r15_7_ ;
  wire  execution_unit_0.register_file_0.r15_8_ ;
  wire  execution_unit_0.register_file_0.r15_9_ ;
  wire  execution_unit_0.register_file_0.r1_10_ ;
  wire  execution_unit_0.register_file_0.r1_11_ ;
  wire  execution_unit_0.register_file_0.r1_12_ ;
  wire  execution_unit_0.register_file_0.r1_13_ ;
  wire  execution_unit_0.register_file_0.r1_14_ ;
  wire  execution_unit_0.register_file_0.r1_15_ ;
  wire  execution_unit_0.register_file_0.r1_1_ ;
  wire  execution_unit_0.register_file_0.r1_2_ ;
  wire  execution_unit_0.register_file_0.r1_3_ ;
  wire  execution_unit_0.register_file_0.r1_4_ ;
  wire  execution_unit_0.register_file_0.r1_5_ ;
  wire  execution_unit_0.register_file_0.r1_6_ ;
  wire  execution_unit_0.register_file_0.r1_7_ ;
  wire  execution_unit_0.register_file_0.r1_8_ ;
  wire  execution_unit_0.register_file_0.r1_9_ ;
  wire  execution_unit_0.register_file_0.r2_4_ ;
  wire  execution_unit_0.register_file_0.r3_0_ ;
  wire  execution_unit_0.register_file_0.r3_10_ ;
  wire  execution_unit_0.register_file_0.r3_11_ ;
  wire  execution_unit_0.register_file_0.r3_12_ ;
  wire  execution_unit_0.register_file_0.r3_13_ ;
  wire  execution_unit_0.register_file_0.r3_14_ ;
  wire  execution_unit_0.register_file_0.r3_15_ ;
  wire  execution_unit_0.register_file_0.r3_1_ ;
  wire  execution_unit_0.register_file_0.r3_2_ ;
  wire  execution_unit_0.register_file_0.r3_3_ ;
  wire  execution_unit_0.register_file_0.r3_4_ ;
  wire  execution_unit_0.register_file_0.r3_5_ ;
  wire  execution_unit_0.register_file_0.r3_6_ ;
  wire  execution_unit_0.register_file_0.r3_7_ ;
  wire  execution_unit_0.register_file_0.r3_8_ ;
  wire  execution_unit_0.register_file_0.r3_9_ ;
  wire  execution_unit_0.register_file_0.r4_0_ ;
  wire  execution_unit_0.register_file_0.r4_10_ ;
  wire  execution_unit_0.register_file_0.r4_11_ ;
  wire  execution_unit_0.register_file_0.r4_12_ ;
  wire  execution_unit_0.register_file_0.r4_13_ ;
  wire  execution_unit_0.register_file_0.r4_14_ ;
  wire  execution_unit_0.register_file_0.r4_15_ ;
  wire  execution_unit_0.register_file_0.r4_1_ ;
  wire  execution_unit_0.register_file_0.r4_2_ ;
  wire  execution_unit_0.register_file_0.r4_3_ ;
  wire  execution_unit_0.register_file_0.r4_4_ ;
  wire  execution_unit_0.register_file_0.r4_5_ ;
  wire  execution_unit_0.register_file_0.r4_6_ ;
  wire  execution_unit_0.register_file_0.r4_7_ ;
  wire  execution_unit_0.register_file_0.r4_8_ ;
  wire  execution_unit_0.register_file_0.r4_9_ ;
  wire  execution_unit_0.register_file_0.r5_0_ ;
  wire  execution_unit_0.register_file_0.r5_10_ ;
  wire  execution_unit_0.register_file_0.r5_11_ ;
  wire  execution_unit_0.register_file_0.r5_12_ ;
  wire  execution_unit_0.register_file_0.r5_13_ ;
  wire  execution_unit_0.register_file_0.r5_14_ ;
  wire  execution_unit_0.register_file_0.r5_15_ ;
  wire  execution_unit_0.register_file_0.r5_1_ ;
  wire  execution_unit_0.register_file_0.r5_2_ ;
  wire  execution_unit_0.register_file_0.r5_3_ ;
  wire  execution_unit_0.register_file_0.r5_4_ ;
  wire  execution_unit_0.register_file_0.r5_5_ ;
  wire  execution_unit_0.register_file_0.r5_6_ ;
  wire  execution_unit_0.register_file_0.r5_7_ ;
  wire  execution_unit_0.register_file_0.r5_8_ ;
  wire  execution_unit_0.register_file_0.r5_9_ ;
  wire  execution_unit_0.register_file_0.r6_0_ ;
  wire  execution_unit_0.register_file_0.r6_10_ ;
  wire  execution_unit_0.register_file_0.r6_11_ ;
  wire  execution_unit_0.register_file_0.r6_12_ ;
  wire  execution_unit_0.register_file_0.r6_13_ ;
  wire  execution_unit_0.register_file_0.r6_14_ ;
  wire  execution_unit_0.register_file_0.r6_15_ ;
  wire  execution_unit_0.register_file_0.r6_1_ ;
  wire  execution_unit_0.register_file_0.r6_2_ ;
  wire  execution_unit_0.register_file_0.r6_3_ ;
  wire  execution_unit_0.register_file_0.r6_4_ ;
  wire  execution_unit_0.register_file_0.r6_5_ ;
  wire  execution_unit_0.register_file_0.r6_6_ ;
  wire  execution_unit_0.register_file_0.r6_7_ ;
  wire  execution_unit_0.register_file_0.r6_8_ ;
  wire  execution_unit_0.register_file_0.r6_9_ ;
  wire  execution_unit_0.register_file_0.r7_0_ ;
  wire  execution_unit_0.register_file_0.r7_10_ ;
  wire  execution_unit_0.register_file_0.r7_11_ ;
  wire  execution_unit_0.register_file_0.r7_12_ ;
  wire  execution_unit_0.register_file_0.r7_13_ ;
  wire  execution_unit_0.register_file_0.r7_14_ ;
  wire  execution_unit_0.register_file_0.r7_15_ ;
  wire  execution_unit_0.register_file_0.r7_1_ ;
  wire  execution_unit_0.register_file_0.r7_2_ ;
  wire  execution_unit_0.register_file_0.r7_3_ ;
  wire  execution_unit_0.register_file_0.r7_4_ ;
  wire  execution_unit_0.register_file_0.r7_5_ ;
  wire  execution_unit_0.register_file_0.r7_6_ ;
  wire  execution_unit_0.register_file_0.r7_7_ ;
  wire  execution_unit_0.register_file_0.r7_8_ ;
  wire  execution_unit_0.register_file_0.r7_9_ ;
  wire  execution_unit_0.register_file_0.r8_0_ ;
  wire  execution_unit_0.register_file_0.r8_10_ ;
  wire  execution_unit_0.register_file_0.r8_11_ ;
  wire  execution_unit_0.register_file_0.r8_12_ ;
  wire  execution_unit_0.register_file_0.r8_13_ ;
  wire  execution_unit_0.register_file_0.r8_14_ ;
  wire  execution_unit_0.register_file_0.r8_15_ ;
  wire  execution_unit_0.register_file_0.r8_1_ ;
  wire  execution_unit_0.register_file_0.r8_2_ ;
  wire  execution_unit_0.register_file_0.r8_3_ ;
  wire  execution_unit_0.register_file_0.r8_4_ ;
  wire  execution_unit_0.register_file_0.r8_5_ ;
  wire  execution_unit_0.register_file_0.r8_6_ ;
  wire  execution_unit_0.register_file_0.r8_7_ ;
  wire  execution_unit_0.register_file_0.r8_8_ ;
  wire  execution_unit_0.register_file_0.r8_9_ ;
  wire  execution_unit_0.register_file_0.r9_0_ ;
  wire  execution_unit_0.register_file_0.r9_10_ ;
  wire  execution_unit_0.register_file_0.r9_11_ ;
  wire  execution_unit_0.register_file_0.r9_12_ ;
  wire  execution_unit_0.register_file_0.r9_13_ ;
  wire  execution_unit_0.register_file_0.r9_14_ ;
  wire  execution_unit_0.register_file_0.r9_15_ ;
  wire  execution_unit_0.register_file_0.r9_1_ ;
  wire  execution_unit_0.register_file_0.r9_2_ ;
  wire  execution_unit_0.register_file_0.r9_3_ ;
  wire  execution_unit_0.register_file_0.r9_4_ ;
  wire  execution_unit_0.register_file_0.r9_5_ ;
  wire  execution_unit_0.register_file_0.r9_6_ ;
  wire  execution_unit_0.register_file_0.r9_7_ ;
  wire  execution_unit_0.register_file_0.r9_8_ ;
  wire  execution_unit_0.register_file_0.r9_9_ ;
  wire  frontend_0.e_state_nxt_0_ ;
  wire  frontend_0.e_state_nxt_1_ ;
  wire  frontend_0.e_state_nxt_2_ ;
  wire  frontend_0.e_state_nxt_3_ ;
  wire  frontend_0.exec_dext_rdy ;
  wire  frontend_0.exec_dst_wr ;
  wire  frontend_0.exec_jmp ;
  wire  frontend_0.exec_src_wr ;
  wire  frontend_0.fe_pmem_wait ;
  wire  frontend_0.i_state_0_ ;
  wire  frontend_0.i_state_1_ ;
  wire  frontend_0.i_state_2_ ;
  wire  frontend_0.i_state_nxt_0_ ;
  wire  frontend_0.i_state_nxt_1_ ;
  wire  frontend_0.i_state_nxt_2_ ;
  wire  frontend_0.inst_dest_bin_0_ ;
  wire  frontend_0.inst_dest_bin_1_ ;
  wire  frontend_0.inst_dest_bin_2_ ;
  wire  frontend_0.inst_dest_bin_3_ ;
  wire  frontend_0.inst_jmp_bin_0_ ;
  wire  frontend_0.inst_jmp_bin_1_ ;
  wire  frontend_0.inst_jmp_bin_2_ ;
  wire  frontend_0.inst_src_bin_0_ ;
  wire  frontend_0.inst_src_bin_1_ ;
  wire  frontend_0.inst_sz_0_ ;
  wire  frontend_0.inst_sz_1_ ;
  wire  frontend_0.irq_addr_1_ ;
  wire  frontend_0.irq_addr_2_ ;
  wire  frontend_0.irq_addr_3_ ;
  wire  frontend_0.irq_addr_4_ ;
  wire  frontend_0.mb_en ;
  wire  frontend_0.pmem_busy ;
  wire  frontend_0.wdt_irq ;
  input irq_0_;
  wire irq_0_;
  input irq_10_;
  wire irq_10_;
  input irq_11_;
  wire irq_11_;
  input irq_12_;
  wire irq_12_;
  input irq_13_;
  wire irq_13_;
  input irq_1_;
  wire irq_1_;
  input irq_2_;
  wire irq_2_;
  input irq_3_;
  wire irq_3_;
  input irq_4_;
  wire irq_4_;
  input irq_5_;
  wire irq_5_;
  input irq_6_;
  wire irq_6_;
  input irq_7_;
  wire irq_7_;
  input irq_8_;
  wire irq_8_;
  input irq_9_;
  wire irq_9_;
  output irq_acc_0_;
  wire irq_acc_0_;
  output irq_acc_10_;
  wire irq_acc_10_;
  output irq_acc_11_;
  wire irq_acc_11_;
  output irq_acc_12_;
  wire irq_acc_12_;
  output irq_acc_13_;
  wire irq_acc_13_;
  output irq_acc_1_;
  wire irq_acc_1_;
  output irq_acc_2_;
  wire irq_acc_2_;
  output irq_acc_3_;
  wire irq_acc_3_;
  output irq_acc_4_;
  wire irq_acc_4_;
  output irq_acc_5_;
  wire irq_acc_5_;
  output irq_acc_6_;
  wire irq_acc_6_;
  output irq_acc_7_;
  wire irq_acc_7_;
  output irq_acc_8_;
  wire irq_acc_8_;
  output irq_acc_9_;
  wire irq_acc_9_;
  input lfxt_clk;
  wire lfxt_clk;
  output lfxt_enable;
  wire lfxt_enable;
  output lfxt_wkup;
  wire lfxt_wkup;
  output mclk;
  wire mclk;
  wire  mem_backbone_0.eu_mdb_in_sel_0_ ;
  wire  mem_backbone_0.eu_mdb_in_sel_1_ ;
  wire  mem_backbone_0.eu_per_en ;
  wire  mem_backbone_0.eu_pmem_en ;
  wire  mem_backbone_0.ext_mem_din_sel ;
  wire  mem_backbone_0.ext_per_en ;
  wire  mem_backbone_0.ext_pmem_en ;
  wire  mem_backbone_0.fe_pmem_en ;
  wire  mem_backbone_0.fe_pmem_en_dly ;
  wire  mem_backbone_0.per_dout_0_ ;
  wire  mem_backbone_0.per_dout_10_ ;
  wire  mem_backbone_0.per_dout_11_ ;
  wire  mem_backbone_0.per_dout_12_ ;
  wire  mem_backbone_0.per_dout_13_ ;
  wire  mem_backbone_0.per_dout_14_ ;
  wire  mem_backbone_0.per_dout_15_ ;
  wire  mem_backbone_0.per_dout_1_ ;
  wire  mem_backbone_0.per_dout_2_ ;
  wire  mem_backbone_0.per_dout_3_ ;
  wire  mem_backbone_0.per_dout_4_ ;
  wire  mem_backbone_0.per_dout_5_ ;
  wire  mem_backbone_0.per_dout_6_ ;
  wire  mem_backbone_0.per_dout_7_ ;
  wire  mem_backbone_0.per_dout_8_ ;
  wire  mem_backbone_0.per_dout_9_ ;
  wire  mem_backbone_0.per_dout_val_0_ ;
  wire  mem_backbone_0.per_dout_val_10_ ;
  wire  mem_backbone_0.per_dout_val_11_ ;
  wire  mem_backbone_0.per_dout_val_12_ ;
  wire  mem_backbone_0.per_dout_val_13_ ;
  wire  mem_backbone_0.per_dout_val_14_ ;
  wire  mem_backbone_0.per_dout_val_15_ ;
  wire  mem_backbone_0.per_dout_val_1_ ;
  wire  mem_backbone_0.per_dout_val_2_ ;
  wire  mem_backbone_0.per_dout_val_3_ ;
  wire  mem_backbone_0.per_dout_val_4_ ;
  wire  mem_backbone_0.per_dout_val_5_ ;
  wire  mem_backbone_0.per_dout_val_6_ ;
  wire  mem_backbone_0.per_dout_val_7_ ;
  wire  mem_backbone_0.per_dout_val_8_ ;
  wire  mem_backbone_0.per_dout_val_9_ ;
  wire  mem_backbone_0.pmem_dout_bckup_0_ ;
  wire  mem_backbone_0.pmem_dout_bckup_10_ ;
  wire  mem_backbone_0.pmem_dout_bckup_11_ ;
  wire  mem_backbone_0.pmem_dout_bckup_12_ ;
  wire  mem_backbone_0.pmem_dout_bckup_13_ ;
  wire  mem_backbone_0.pmem_dout_bckup_14_ ;
  wire  mem_backbone_0.pmem_dout_bckup_15_ ;
  wire  mem_backbone_0.pmem_dout_bckup_1_ ;
  wire  mem_backbone_0.pmem_dout_bckup_2_ ;
  wire  mem_backbone_0.pmem_dout_bckup_3_ ;
  wire  mem_backbone_0.pmem_dout_bckup_4_ ;
  wire  mem_backbone_0.pmem_dout_bckup_5_ ;
  wire  mem_backbone_0.pmem_dout_bckup_6_ ;
  wire  mem_backbone_0.pmem_dout_bckup_7_ ;
  wire  mem_backbone_0.pmem_dout_bckup_8_ ;
  wire  mem_backbone_0.pmem_dout_bckup_9_ ;
  wire  mem_backbone_0.pmem_dout_bckup_sel ;
  wire  multiplier_0.acc_sel ;
  wire  multiplier_0.cycle_0_ ;
  wire  multiplier_0.cycle_1_ ;
  wire  multiplier_0.op1_0_ ;
  wire  multiplier_0.op1_10_ ;
  wire  multiplier_0.op1_11_ ;
  wire  multiplier_0.op1_12_ ;
  wire  multiplier_0.op1_13_ ;
  wire  multiplier_0.op1_14_ ;
  wire  multiplier_0.op1_15_ ;
  wire  multiplier_0.op1_1_ ;
  wire  multiplier_0.op1_2_ ;
  wire  multiplier_0.op1_3_ ;
  wire  multiplier_0.op1_4_ ;
  wire  multiplier_0.op1_5_ ;
  wire  multiplier_0.op1_6_ ;
  wire  multiplier_0.op1_7_ ;
  wire  multiplier_0.op1_8_ ;
  wire  multiplier_0.op1_9_ ;
  wire  multiplier_0.op2_0_ ;
  wire  multiplier_0.op2_10_ ;
  wire  multiplier_0.op2_11_ ;
  wire  multiplier_0.op2_12_ ;
  wire  multiplier_0.op2_13_ ;
  wire  multiplier_0.op2_14_ ;
  wire  multiplier_0.op2_15_ ;
  wire  multiplier_0.op2_1_ ;
  wire  multiplier_0.op2_2_ ;
  wire  multiplier_0.op2_3_ ;
  wire  multiplier_0.op2_4_ ;
  wire  multiplier_0.op2_5_ ;
  wire  multiplier_0.op2_6_ ;
  wire  multiplier_0.op2_7_ ;
  wire  multiplier_0.op2_8_ ;
  wire  multiplier_0.op2_9_ ;
  wire  multiplier_0.op2_wr ;
  wire  multiplier_0.per_dout_0_ ;
  wire  multiplier_0.per_dout_10_ ;
  wire  multiplier_0.per_dout_11_ ;
  wire  multiplier_0.per_dout_12_ ;
  wire  multiplier_0.per_dout_13_ ;
  wire  multiplier_0.per_dout_14_ ;
  wire  multiplier_0.per_dout_15_ ;
  wire  multiplier_0.per_dout_1_ ;
  wire  multiplier_0.per_dout_2_ ;
  wire  multiplier_0.per_dout_3_ ;
  wire  multiplier_0.per_dout_4_ ;
  wire  multiplier_0.per_dout_5_ ;
  wire  multiplier_0.per_dout_6_ ;
  wire  multiplier_0.per_dout_7_ ;
  wire  multiplier_0.per_dout_8_ ;
  wire  multiplier_0.per_dout_9_ ;
  wire  multiplier_0.reshi_0_ ;
  wire  multiplier_0.reshi_10_ ;
  wire  multiplier_0.reshi_11_ ;
  wire  multiplier_0.reshi_12_ ;
  wire  multiplier_0.reshi_13_ ;
  wire  multiplier_0.reshi_14_ ;
  wire  multiplier_0.reshi_15_ ;
  wire  multiplier_0.reshi_1_ ;
  wire  multiplier_0.reshi_2_ ;
  wire  multiplier_0.reshi_3_ ;
  wire  multiplier_0.reshi_4_ ;
  wire  multiplier_0.reshi_5_ ;
  wire  multiplier_0.reshi_6_ ;
  wire  multiplier_0.reshi_7_ ;
  wire  multiplier_0.reshi_8_ ;
  wire  multiplier_0.reshi_9_ ;
  wire  multiplier_0.reslo_0_ ;
  wire  multiplier_0.reslo_10_ ;
  wire  multiplier_0.reslo_11_ ;
  wire  multiplier_0.reslo_12_ ;
  wire  multiplier_0.reslo_13_ ;
  wire  multiplier_0.reslo_14_ ;
  wire  multiplier_0.reslo_15_ ;
  wire  multiplier_0.reslo_1_ ;
  wire  multiplier_0.reslo_2_ ;
  wire  multiplier_0.reslo_3_ ;
  wire  multiplier_0.reslo_4_ ;
  wire  multiplier_0.reslo_5_ ;
  wire  multiplier_0.reslo_6_ ;
  wire  multiplier_0.reslo_7_ ;
  wire  multiplier_0.reslo_8_ ;
  wire  multiplier_0.reslo_9_ ;
  wire  multiplier_0.sign_sel ;
  wire  multiplier_0.sumext_0_ ;
  wire  multiplier_0.sumext_10_ ;
  input nmi;
  wire nmi;
  output per_addr_0_;
  wire per_addr_0_;
  output per_addr_10_;
  wire per_addr_10_;
  output per_addr_11_;
  wire per_addr_11_;
  output per_addr_12_;
  wire per_addr_12_;
  output per_addr_13_;
  wire per_addr_13_;
  output per_addr_1_;
  wire per_addr_1_;
  output per_addr_2_;
  wire per_addr_2_;
  output per_addr_3_;
  wire per_addr_3_;
  output per_addr_4_;
  wire per_addr_4_;
  output per_addr_5_;
  wire per_addr_5_;
  output per_addr_6_;
  wire per_addr_6_;
  output per_addr_7_;
  wire per_addr_7_;
  output per_addr_8_;
  wire per_addr_8_;
  output per_addr_9_;
  wire per_addr_9_;
  output per_din_0_;
  wire per_din_0_;
  output per_din_10_;
  wire per_din_10_;
  output per_din_11_;
  wire per_din_11_;
  output per_din_12_;
  wire per_din_12_;
  output per_din_13_;
  wire per_din_13_;
  output per_din_14_;
  wire per_din_14_;
  output per_din_15_;
  wire per_din_15_;
  output per_din_1_;
  wire per_din_1_;
  output per_din_2_;
  wire per_din_2_;
  output per_din_3_;
  wire per_din_3_;
  output per_din_4_;
  wire per_din_4_;
  output per_din_5_;
  wire per_din_5_;
  output per_din_6_;
  wire per_din_6_;
  output per_din_7_;
  wire per_din_7_;
  output per_din_8_;
  wire per_din_8_;
  output per_din_9_;
  wire per_din_9_;
  input per_dout_0_;
  wire per_dout_0_;
  input per_dout_10_;
  wire per_dout_10_;
  input per_dout_11_;
  wire per_dout_11_;
  input per_dout_12_;
  wire per_dout_12_;
  input per_dout_13_;
  wire per_dout_13_;
  input per_dout_14_;
  wire per_dout_14_;
  input per_dout_15_;
  wire per_dout_15_;
  input per_dout_1_;
  wire per_dout_1_;
  input per_dout_2_;
  wire per_dout_2_;
  input per_dout_3_;
  wire per_dout_3_;
  input per_dout_4_;
  wire per_dout_4_;
  input per_dout_5_;
  wire per_dout_5_;
  input per_dout_6_;
  wire per_dout_6_;
  input per_dout_7_;
  wire per_dout_7_;
  input per_dout_8_;
  wire per_dout_8_;
  input per_dout_9_;
  wire per_dout_9_;
  output per_en;
  wire per_en;
  output per_we_0_;
  wire per_we_0_;
  output per_we_1_;
  wire per_we_1_;
  output pmem_addr_0_;
  wire pmem_addr_0_;
  output pmem_addr_10_;
  wire pmem_addr_10_;
  output pmem_addr_11_;
  wire pmem_addr_11_;
  output pmem_addr_12_;
  wire pmem_addr_12_;
  output pmem_addr_13_;
  wire pmem_addr_13_;
  output pmem_addr_1_;
  wire pmem_addr_1_;
  output pmem_addr_2_;
  wire pmem_addr_2_;
  output pmem_addr_3_;
  wire pmem_addr_3_;
  output pmem_addr_4_;
  wire pmem_addr_4_;
  output pmem_addr_5_;
  wire pmem_addr_5_;
  output pmem_addr_6_;
  wire pmem_addr_6_;
  output pmem_addr_7_;
  wire pmem_addr_7_;
  output pmem_addr_8_;
  wire pmem_addr_8_;
  output pmem_addr_9_;
  wire pmem_addr_9_;
  output pmem_cen;
  wire pmem_cen;
  output pmem_din_0_;
  wire pmem_din_0_;
  output pmem_din_10_;
  wire pmem_din_10_;
  output pmem_din_11_;
  wire pmem_din_11_;
  output pmem_din_12_;
  wire pmem_din_12_;
  output pmem_din_13_;
  wire pmem_din_13_;
  output pmem_din_14_;
  wire pmem_din_14_;
  output pmem_din_15_;
  wire pmem_din_15_;
  output pmem_din_1_;
  wire pmem_din_1_;
  output pmem_din_2_;
  wire pmem_din_2_;
  output pmem_din_3_;
  wire pmem_din_3_;
  output pmem_din_4_;
  wire pmem_din_4_;
  output pmem_din_5_;
  wire pmem_din_5_;
  output pmem_din_6_;
  wire pmem_din_6_;
  output pmem_din_7_;
  wire pmem_din_7_;
  output pmem_din_8_;
  wire pmem_din_8_;
  output pmem_din_9_;
  wire pmem_din_9_;
  input pmem_dout_0_;
  wire pmem_dout_0_;
  input pmem_dout_10_;
  wire pmem_dout_10_;
  input pmem_dout_11_;
  wire pmem_dout_11_;
  input pmem_dout_12_;
  wire pmem_dout_12_;
  input pmem_dout_13_;
  wire pmem_dout_13_;
  input pmem_dout_14_;
  wire pmem_dout_14_;
  input pmem_dout_15_;
  wire pmem_dout_15_;
  input pmem_dout_1_;
  wire pmem_dout_1_;
  input pmem_dout_2_;
  wire pmem_dout_2_;
  input pmem_dout_3_;
  wire pmem_dout_3_;
  input pmem_dout_4_;
  wire pmem_dout_4_;
  input pmem_dout_5_;
  wire pmem_dout_5_;
  input pmem_dout_6_;
  wire pmem_dout_6_;
  input pmem_dout_7_;
  wire pmem_dout_7_;
  input pmem_dout_8_;
  wire pmem_dout_8_;
  input pmem_dout_9_;
  wire pmem_dout_9_;
  output pmem_wen_0_;
  wire pmem_wen_0_;
  output pmem_wen_1_;
  wire pmem_wen_1_;
  output puc_rst;
  wire puc_rst;
  input reset_n;
  wire reset_n;
  input scan_enable;
  wire scan_enable;
  input scan_mode;
  wire scan_mode;
  wire  sfr_0.cpu_nr_rd_10_ ;
  wire  sfr_0.cpu_nr_rd_11_ ;
  wire  sfr_0.cpu_nr_rd_12_ ;
  wire  sfr_0.cpu_nr_rd_13_ ;
  wire  sfr_0.cpu_nr_rd_2_ ;
  wire  sfr_0.cpu_nr_rd_3_ ;
  wire  sfr_0.cpu_nr_rd_4_ ;
  wire  sfr_0.cpu_nr_rd_5_ ;
  wire  sfr_0.cpu_nr_rd_6_ ;
  wire  sfr_0.cpu_nr_rd_7_ ;
  wire  sfr_0.cpu_nr_rd_9_ ;
  wire  sfr_0.ie1_0_ ;
  wire  sfr_0.ifg1_0_ ;
  wire  sfr_0.per_dout_0_ ;
  wire  sfr_0.per_dout_14_ ;
  wire  sfr_0.per_dout_15_ ;
  wire  sfr_0.per_dout_1_ ;
  wire  sfr_0.per_dout_8_ ;
  wire  sfr_0.wdtifg_sw_clr ;
  wire  sfr_0.wdtifg_sw_set ;
  output smclk;
  wire smclk;
  output smclk_en;
  wire smclk_en;
  wire  watchdog_0.per_dout_0_ ;
  wire  watchdog_0.per_dout_11_ ;
  wire  watchdog_0.per_dout_1_ ;
  wire  watchdog_0.per_dout_2_ ;
  wire  watchdog_0.per_dout_4_ ;
  wire  watchdog_0.per_dout_7_ ;
  wire  watchdog_0.wdtcnt_0_ ;
  wire  watchdog_0.wdtcnt_10_ ;
  wire  watchdog_0.wdtcnt_11_ ;
  wire  watchdog_0.wdtcnt_12_ ;
  wire  watchdog_0.wdtcnt_13_ ;
  wire  watchdog_0.wdtcnt_14_ ;
  wire  watchdog_0.wdtcnt_15_ ;
  wire  watchdog_0.wdtcnt_1_ ;
  wire  watchdog_0.wdtcnt_2_ ;
  wire  watchdog_0.wdtcnt_3_ ;
  wire  watchdog_0.wdtcnt_4_ ;
  wire  watchdog_0.wdtcnt_5_ ;
  wire  watchdog_0.wdtcnt_6_ ;
  wire  watchdog_0.wdtcnt_7_ ;
  wire  watchdog_0.wdtcnt_8_ ;
  wire  watchdog_0.wdtcnt_9_ ;
  wire  watchdog_0.wdtctl_0_ ;
  wire  watchdog_0.wdtctl_1_ ;
  wire  watchdog_0.wdtctl_2_ ;
  wire  watchdog_0.wdtctl_4_ ;
  wire  watchdog_0.wdtctl_7_ ;
  input wkup;
  wire wkup;
  INVX1 _06329_ (
    .A( multiplier_0.per_dout_0_ ),
    .Y(_00045_)
  );
  INVX1 _06330_ (
    .A( multiplier_0.per_dout_1_ ),
    .Y(_00046_)
  );
  INVX1 _06331_ (
    .A( multiplier_0.per_dout_2_ ),
    .Y(_00047_)
  );
  INVX1 _06332_ (
    .A( multiplier_0.per_dout_3_ ),
    .Y(_00000_)
  );
  INVX1 _06333_ (
    .A( multiplier_0.per_dout_4_ ),
    .Y(_00001_)
  );
  INVX1 _06334_ (
    .A( multiplier_0.per_dout_5_ ),
    .Y(_00002_)
  );
  INVX1 _06335_ (
    .A( multiplier_0.per_dout_6_ ),
    .Y(_00003_)
  );
  INVX1 _06336_ (
    .A( multiplier_0.per_dout_7_ ),
    .Y(_00004_)
  );
  INVX1 _06337_ (
    .A( multiplier_0.per_dout_8_ ),
    .Y(_00005_)
  );
  INVX1 _06338_ (
    .A( multiplier_0.per_dout_9_ ),
    .Y(_00006_)
  );
  INVX1 _06339_ (
    .A( multiplier_0.per_dout_10_ ),
    .Y(_00007_)
  );
  INVX1 _06340_ (
    .A( multiplier_0.per_dout_11_ ),
    .Y(_00008_)
  );
  INVX1 _06341_ (
    .A( multiplier_0.per_dout_12_ ),
    .Y(_00009_)
  );
  INVX1 _06342_ (
    .A( multiplier_0.per_dout_13_ ),
    .Y(_00010_)
  );
  INVX1 _06343_ (
    .A( multiplier_0.per_dout_14_ ),
    .Y(_00011_)
  );
  INVX1 _06344_ (
    .A( multiplier_0.per_dout_15_ ),
    .Y(_00012_)
  );
  NOR2X1 _06345_ (
    .A(1'h0),
    .B(per_dout_0_),
    .Y(_00013_)
  );
  NOR2X1 _06346_ (
    .A( sfr_0.per_dout_0_ ),
    .B( watchdog_0.per_dout_0_ ),
    .Y(_00014_)
  );
  NAND3X1 _06347_ (
    .A(_00045_),
    .B(_00013_),
    .C(_00014_),
    .Y( mem_backbone_0.per_dout_0_ )
  );
  NOR2X1 _06348_ (
    .A( clock_module_0.bcsctl2_rd_1_ ),
    .B(per_dout_1_),
    .Y(_00015_)
  );
  NOR2X1 _06349_ (
    .A( sfr_0.per_dout_1_ ),
    .B( watchdog_0.per_dout_1_ ),
    .Y(_00016_)
  );
  NAND3X1 _06350_ (
    .A(_00046_),
    .B(_00015_),
    .C(_00016_),
    .Y( mem_backbone_0.per_dout_1_ )
  );
  NOR2X1 _06351_ (
    .A( clock_module_0.bcsctl2_rd_2_ ),
    .B(per_dout_2_),
    .Y(_00017_)
  );
  NOR2X1 _06352_ (
    .A( sfr_0.cpu_nr_rd_2_ ),
    .B( watchdog_0.per_dout_2_ ),
    .Y(_00018_)
  );
  NAND3X1 _06353_ (
    .A(_00047_),
    .B(_00017_),
    .C(_00018_),
    .Y( mem_backbone_0.per_dout_2_ )
  );
  NOR2X1 _06354_ (
    .A( clock_module_0.bcsctl2_rd_3_ ),
    .B(per_dout_3_),
    .Y(_00019_)
  );
  NOR2X1 _06355_ (
    .A( sfr_0.cpu_nr_rd_3_ ),
    .B(1'h0),
    .Y(_00020_)
  );
  NAND3X1 _06356_ (
    .A(_00000_),
    .B(_00019_),
    .C(_00020_),
    .Y( mem_backbone_0.per_dout_3_ )
  );
  NOR2X1 _06357_ (
    .A(1'h0),
    .B(per_dout_4_),
    .Y(_00021_)
  );
  NOR2X1 _06358_ (
    .A( sfr_0.cpu_nr_rd_4_ ),
    .B( watchdog_0.per_dout_4_ ),
    .Y(_00022_)
  );
  NAND3X1 _06359_ (
    .A(_00001_),
    .B(_00021_),
    .C(_00022_),
    .Y( mem_backbone_0.per_dout_4_ )
  );
  NOR2X1 _06360_ (
    .A(1'h0),
    .B(per_dout_5_),
    .Y(_00023_)
  );
  NOR2X1 _06361_ (
    .A( sfr_0.cpu_nr_rd_5_ ),
    .B(1'h0),
    .Y(_00024_)
  );
  NAND3X1 _06362_ (
    .A(_00002_),
    .B(_00023_),
    .C(_00024_),
    .Y( mem_backbone_0.per_dout_5_ )
  );
  NOR2X1 _06363_ (
    .A(1'h0),
    .B(per_dout_6_),
    .Y(_00025_)
  );
  NOR2X1 _06364_ (
    .A( sfr_0.cpu_nr_rd_6_ ),
    .B(1'h0),
    .Y(_00026_)
  );
  NAND3X1 _06365_ (
    .A(_00003_),
    .B(_00025_),
    .C(_00026_),
    .Y( mem_backbone_0.per_dout_6_ )
  );
  NOR2X1 _06366_ (
    .A(1'h0),
    .B(per_dout_7_),
    .Y(_00027_)
  );
  NOR2X1 _06367_ (
    .A( sfr_0.cpu_nr_rd_7_ ),
    .B( watchdog_0.per_dout_7_ ),
    .Y(_00028_)
  );
  NAND3X1 _06368_ (
    .A(_00004_),
    .B(_00027_),
    .C(_00028_),
    .Y( mem_backbone_0.per_dout_7_ )
  );
  NOR2X1 _06369_ (
    .A(1'h0),
    .B(per_dout_8_),
    .Y(_00029_)
  );
  NOR2X1 _06370_ (
    .A( sfr_0.per_dout_8_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00030_)
  );
  NAND3X1 _06371_ (
    .A(_00005_),
    .B(_00029_),
    .C(_00030_),
    .Y( mem_backbone_0.per_dout_8_ )
  );
  NOR2X1 _06372_ (
    .A(1'h0),
    .B(per_dout_9_),
    .Y(_00031_)
  );
  NOR2X1 _06373_ (
    .A( sfr_0.cpu_nr_rd_9_ ),
    .B(1'h0),
    .Y(_00032_)
  );
  NAND3X1 _06374_ (
    .A(_00006_),
    .B(_00031_),
    .C(_00032_),
    .Y( mem_backbone_0.per_dout_9_ )
  );
  NOR2X1 _06375_ (
    .A(1'h0),
    .B(per_dout_10_),
    .Y(_00033_)
  );
  NOR2X1 _06376_ (
    .A( sfr_0.cpu_nr_rd_10_ ),
    .B(1'h0),
    .Y(_00034_)
  );
  NAND3X1 _06377_ (
    .A(_00007_),
    .B(_00033_),
    .C(_00034_),
    .Y( mem_backbone_0.per_dout_10_ )
  );
  NOR2X1 _06378_ (
    .A(1'h0),
    .B(per_dout_11_),
    .Y(_00035_)
  );
  NOR2X1 _06379_ (
    .A( sfr_0.cpu_nr_rd_11_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00036_)
  );
  NAND3X1 _06380_ (
    .A(_00008_),
    .B(_00035_),
    .C(_00036_),
    .Y( mem_backbone_0.per_dout_11_ )
  );
  NOR2X1 _06381_ (
    .A( clock_module_0.bcsctl1_rd_12_ ),
    .B(per_dout_12_),
    .Y(_00037_)
  );
  NOR2X1 _06382_ (
    .A( sfr_0.cpu_nr_rd_12_ ),
    .B(1'h0),
    .Y(_00038_)
  );
  NAND3X1 _06383_ (
    .A(_00009_),
    .B(_00037_),
    .C(_00038_),
    .Y( mem_backbone_0.per_dout_12_ )
  );
  NOR2X1 _06384_ (
    .A( clock_module_0.bcsctl1_rd_13_ ),
    .B(per_dout_13_),
    .Y(_00039_)
  );
  NOR2X1 _06385_ (
    .A( sfr_0.cpu_nr_rd_13_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00040_)
  );
  NAND3X1 _06386_ (
    .A(_00010_),
    .B(_00039_),
    .C(_00040_),
    .Y( mem_backbone_0.per_dout_13_ )
  );
  NOR2X1 _06387_ (
    .A(1'h0),
    .B(per_dout_14_),
    .Y(_00041_)
  );
  NOR2X1 _06388_ (
    .A( sfr_0.per_dout_14_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00042_)
  );
  NAND3X1 _06389_ (
    .A(_00011_),
    .B(_00041_),
    .C(_00042_),
    .Y( mem_backbone_0.per_dout_14_ )
  );
  NOR2X1 _06390_ (
    .A(1'h0),
    .B(per_dout_15_),
    .Y(_00043_)
  );
  NOR2X1 _06391_ (
    .A( sfr_0.per_dout_15_ ),
    .B(1'h0),
    .Y(_00044_)
  );
  NAND3X1 _06392_ (
    .A(_00012_),
    .B(_00043_),
    .C(_00044_),
    .Y( mem_backbone_0.per_dout_15_ )
  );
  INVX1 _06393_ (
    .A( clock_module_0.aclk_div_0_ ),
    .Y(_00099_)
  );
  INVX1 _06394_ (
    .A(reset_n),
    .Y( clock_module_0.por_a )
  );
  INVX1 _06395_ (
    .A(dbg_en),
    .Y( clock_module_0.dbg_rst_nxt )
  );
  INVX1 _06396_ (
    .A( clock_module_0.puc_noscan_n ),
    .Y(_06327_)
  );
  INVX1 _06397_ (
    .A(_06269_),
    .Y(_00100_)
  );
  INVX1 _06398_ (
    .A(_06271_),
    .Y(_00101_)
  );
  INVX1 _06399_ (
    .A(_06265_),
    .Y(_00102_)
  );
  INVX1 _06400_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .Y(_00103_)
  );
  INVX1 _06401_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .Y(_00104_)
  );
  INVX1 _06402_ (
    .A( clock_module_0.lfxt_clk_dly ),
    .Y(_00105_)
  );
  INVX1 _06403_ (
    .A( clock_module_0.oscoff ),
    .Y(_00106_)
  );
  INVX1 _06404_ (
    .A( clock_module_0.aclk_div_1_ ),
    .Y(_00107_)
  );
  INVX1 _06405_ (
    .A( clock_module_0.smclk_div_1_ ),
    .Y(_00108_)
  );
  INVX1 _06406_ (
    .A( clock_module_0.smclk_div_2_ ),
    .Y(_00109_)
  );
  INVX1 _06407_ (
    .A( clock_module_0.por ),
    .Y(_00050_)
  );
  NOR2X1 _06408_ (
    .A( clock_module_0.dbg_rst_nxt ),
    .B( clock_module_0.puc_noscan_n ),
    .Y(_00110_)
  );
  AOI21X1 _06409_ (
    .A( clock_module_0.dbg_rst ),
    .B(_00110_),
    .C( clock_module_0.dbg_cpu_reset ),
    .Y( clock_module_0.sync_cell_puc.data_in )
  );
  NOR2X1 _06410_ (
    .A(_06264_),
    .B(1'h0),
    .Y(_00111_)
  );
  NAND3X1 _06411_ (
    .A(_00102_),
    .B(_06291_),
    .C(_00111_),
    .Y(_00112_)
  );
  INVX1 _06412_ (
    .A(_00112_),
    .Y(_00113_)
  );
  NOR2X1 _06413_ (
    .A(_06273_),
    .B(_06272_),
    .Y(_00114_)
  );
  NOR2X1 _06414_ (
    .A(_06263_),
    .B(_06274_),
    .Y(_00115_)
  );
  NAND2X1 _06415_ (
    .A(_00114_),
    .B(_00115_),
    .Y(_00116_)
  );
  NAND2X1 _06416_ (
    .A(_00100_),
    .B(_06268_),
    .Y(_00117_)
  );
  NAND2X1 _06417_ (
    .A(_00101_),
    .B(_06270_),
    .Y(_00118_)
  );
  NOR3X1 _06418_ (
    .A(_00116_),
    .B(_00117_),
    .C(_00118_),
    .Y(_00119_)
  );
  NOR2X1 _06419_ (
    .A(_06293_),
    .B(_06292_),
    .Y(_00120_)
  );
  NAND3X1 _06420_ (
    .A(_00113_),
    .B(_00119_),
    .C(_00120_),
    .Y(_00121_)
  );
  NOR2X1 _06421_ (
    .A(_06266_),
    .B(_06262_),
    .Y(_00122_)
  );
  AND2X1 _06422_ (
    .A(_06267_),
    .B(_00122_),
    .Y(_00063_)
  );
  NAND2X1 _06423_ (
    .A(_06267_),
    .B(_00122_),
    .Y(_00064_)
  );
  NOR2X1 _06424_ (
    .A(_00121_),
    .B(_00064_),
    .Y(_00065_)
  );
  AND2X1 _06425_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_00065_),
    .Y( clock_module_0.bcsctl2_rd_1_ )
  );
  AND2X1 _06426_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .B(_00065_),
    .Y( clock_module_0.bcsctl2_rd_2_ )
  );
  AND2X1 _06427_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_00065_),
    .Y( clock_module_0.bcsctl2_rd_3_ )
  );
  NAND2X1 _06428_ (
    .A(_06266_),
    .B(_06262_),
    .Y(_00066_)
  );
  NOR2X1 _06429_ (
    .A(_06267_),
    .B(_00066_),
    .Y(_00067_)
  );
  NOR3X1 _06430_ (
    .A(_06267_),
    .B(_00121_),
    .C(_00066_),
    .Y(_00068_)
  );
  AND2X1 _06431_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B(_00068_),
    .Y( clock_module_0.bcsctl1_rd_12_ )
  );
  AND2X1 _06432_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_00068_),
    .Y( clock_module_0.bcsctl1_rd_13_ )
  );
  OAI21X1 _06433_ (
    .A(_00104_),
    .B( clock_module_0.aclk_div_2_ ),
    .C( clock_module_0.aclk_div_1_ ),
    .Y(_00069_)
  );
  OR2X1 _06434_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .Y(_00070_)
  );
  OAI21X1 _06435_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .C(_00099_),
    .Y(_00071_)
  );
  NAND2X1 _06436_ (
    .A(_00105_),
    .B( clock_module_0.lfxt_clk_s ),
    .Y(_00072_)
  );
  NOR2X1 _06437_ (
    .A( clock_module_0.oscoff ),
    .B(_00072_),
    .Y(_00073_)
  );
  NAND3X1 _06438_ (
    .A(_00105_),
    .B( clock_module_0.lfxt_clk_s ),
    .C(_00106_),
    .Y(_00074_)
  );
  NAND3X1 _06439_ (
    .A(cpu_en),
    .B(_00071_),
    .C(_00073_),
    .Y(_00075_)
  );
  AOI21X1 _06440_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_00069_),
    .C(_00075_),
    .Y(_00048_)
  );
  AOI21X1 _06441_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_00074_),
    .C( clock_module_0.scg1 ),
    .Y(_00076_)
  );
  AOI21X1 _06442_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_00109_),
    .C(_00108_),
    .Y(_00077_)
  );
  OR2X1 _06443_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B( clock_module_0.bcsctl2_2_ ),
    .Y(_00078_)
  );
  OAI21X1 _06444_ (
    .A(_00103_),
    .B(_00077_),
    .C( clock_module_0.smclk_div_0_ ),
    .Y(_00079_)
  );
  NAND2X1 _06445_ (
    .A(cpu_en),
    .B(_00076_),
    .Y(_00080_)
  );
  AOI21X1 _06446_ (
    .A(_00078_),
    .B(_00079_),
    .C(_00080_),
    .Y(_00049_)
  );
  OR2X1 _06447_ (
    .A( clock_module_0.wdt_reset ),
    .B( clock_module_0.por ),
    .Y( clock_module_0.puc_a )
  );
  NOR2X1 _06448_ (
    .A(_06273_),
    .B(_06274_),
    .Y(_00081_)
  );
  NAND3X1 _06449_ (
    .A(_00100_),
    .B(_00101_),
    .C(_00081_),
    .Y(_00082_)
  );
  NOR2X1 _06450_ (
    .A(_06272_),
    .B(_06263_),
    .Y(_00083_)
  );
  NAND3X1 _06451_ (
    .A(_06268_),
    .B(_06270_),
    .C(_00083_),
    .Y(_00084_)
  );
  NOR3X1 _06452_ (
    .A(_00112_),
    .B(_00082_),
    .C(_00084_),
    .Y(_00085_)
  );
  NAND3X1 _06453_ (
    .A(_06292_),
    .B(_00063_),
    .C(_00085_),
    .Y(_00086_)
  );
  MUX2X1 _06454_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_06282_),
    .S(_00086_),
    .Y(_00087_)
  );
  INVX1 _06455_ (
    .A(_00087_),
    .Y(_00052_)
  );
  MUX2X1 _06456_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .B(_06283_),
    .S(_00086_),
    .Y(_00088_)
  );
  INVX1 _06457_ (
    .A(_00088_),
    .Y(_00053_)
  );
  MUX2X1 _06458_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_06284_),
    .S(_00086_),
    .Y(_00089_)
  );
  INVX1 _06459_ (
    .A(_00089_),
    .Y(_00054_)
  );
  OAI21X1 _06460_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B( clock_module_0.bcsctl2_2_ ),
    .C(_00076_),
    .Y(_00090_)
  );
  NAND3X1 _06461_ (
    .A( clock_module_0.smclk_div_0_ ),
    .B(_00076_),
    .C(_00078_),
    .Y(_00091_)
  );
  XNOR2X1 _06462_ (
    .A( clock_module_0.smclk_div_0_ ),
    .B(_00090_),
    .Y(_00055_)
  );
  NOR2X1 _06463_ (
    .A(_00108_),
    .B(_00091_),
    .Y(_00092_)
  );
  XNOR2X1 _06464_ (
    .A( clock_module_0.smclk_div_1_ ),
    .B(_00091_),
    .Y(_00056_)
  );
  XNOR2X1 _06465_ (
    .A(_00109_),
    .B(_00092_),
    .Y(_00057_)
  );
  OAI21X1 _06466_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .C(_00073_),
    .Y(_00093_)
  );
  NAND3X1 _06467_ (
    .A( clock_module_0.aclk_div_0_ ),
    .B(_00070_),
    .C(_00073_),
    .Y(_00094_)
  );
  XNOR2X1 _06468_ (
    .A( clock_module_0.aclk_div_0_ ),
    .B(_00093_),
    .Y(_00058_)
  );
  NOR2X1 _06469_ (
    .A(_00107_),
    .B(_00094_),
    .Y(_00095_)
  );
  XNOR2X1 _06470_ (
    .A( clock_module_0.aclk_div_1_ ),
    .B(_00094_),
    .Y(_00059_)
  );
  XOR2X1 _06471_ (
    .A( clock_module_0.aclk_div_2_ ),
    .B(_00095_),
    .Y(_00060_)
  );
  NAND3X1 _06472_ (
    .A(_06293_),
    .B(_00067_),
    .C(_00085_),
    .Y(_00096_)
  );
  MUX2X1 _06473_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B(_06278_),
    .S(_00096_),
    .Y(_00097_)
  );
  INVX1 _06474_ (
    .A(_00097_),
    .Y(_00061_)
  );
  MUX2X1 _06475_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_06279_),
    .S(_00096_),
    .Y(_00098_)
  );
  INVX1 _06476_ (
    .A(_00098_),
    .Y(_00062_)
  );
  INVX1 _06477_ (
    .A( clock_module_0.por ),
    .Y(_00051_)
  );
  DFFSR _06478_ (
    .CLK(dco_clk),
    .D( clock_module_0.dbg_rst_nxt ),
    .Q( clock_module_0.dbg_rst ),
    .R(1'h1),
    .S(_00050_)
  );
  DFFSR _06479_ (
    .CLK(dco_clk),
    .D(_00052_),
    .Q( clock_module_0.bcsctl2_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06480_ (
    .CLK(dco_clk),
    .D(_00053_),
    .Q( clock_module_0.bcsctl2_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06481_ (
    .CLK(dco_clk),
    .D(_00054_),
    .Q( clock_module_0.bcsctl2_3_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06482_ (
    .CLK(dco_clk),
    .D(_00049_),
    .Q(_06328_),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06483_ (
    .CLK(dco_clk),
    .D(_00048_),
    .Q(_06213_),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06484_ (
    .CLK(dco_clk),
    .D(_00055_),
    .Q( clock_module_0.smclk_div_0_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06485_ (
    .CLK(dco_clk),
    .D(_00056_),
    .Q( clock_module_0.smclk_div_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06486_ (
    .CLK(dco_clk),
    .D(_00057_),
    .Q( clock_module_0.smclk_div_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06487_ (
    .CLK(dco_clk),
    .D( clock_module_0.lfxt_clk_s ),
    .Q( clock_module_0.lfxt_clk_dly ),
    .R(_00051_),
    .S(1'h1)
  );
  DFFSR _06488_ (
    .CLK(dco_clk),
    .D(_00058_),
    .Q( clock_module_0.aclk_div_0_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06489_ (
    .CLK(dco_clk),
    .D(_00059_),
    .Q( clock_module_0.aclk_div_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06490_ (
    .CLK(dco_clk),
    .D(_00060_),
    .Q( clock_module_0.aclk_div_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06491_ (
    .CLK(dco_clk),
    .D(_00061_),
    .Q( clock_module_0.bcsctl1_4_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06492_ (
    .CLK(dco_clk),
    .D(_00062_),
    .Q( clock_module_0.bcsctl1_5_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  INVX1 _06493_ (
    .A( clock_module_0.por ),
    .Y(_00123_)
  );
  INVX1 _06494_ (
    .A( clock_module_0.por ),
    .Y(_00124_)
  );
  DFFSR _06495_ (
    .CLK(dco_clk),
    .D(lfxt_clk),
    .Q( clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .R(_00123_),
    .S(1'h1)
  );
  DFFSR _06496_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .Q( clock_module_0.lfxt_clk_s ),
    .R(_00124_),
    .S(1'h1)
  );
  INVX1 _06497_ (
    .A( clock_module_0.puc_a ),
    .Y(_00125_)
  );
  INVX1 _06498_ (
    .A( clock_module_0.puc_a ),
    .Y(_00126_)
  );
  DFFSR _06499_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_puc.data_in ),
    .Q( clock_module_0.sync_cell_puc.data_sync_0_ ),
    .R(_00125_),
    .S(1'h1)
  );
  DFFSR _06500_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_puc.data_sync_0_ ),
    .Q( clock_module_0.puc_noscan_n ),
    .R(_00126_),
    .S(1'h1)
  );
  INVX1 _06501_ (
    .A( clock_module_0.por_a ),
    .Y(_00127_)
  );
  INVX1 _06502_ (
    .A( clock_module_0.por_a ),
    .Y(_00128_)
  );
  DFFSR _06503_ (
    .CLK(dco_clk),
    .D(1'h0),
    .Q( clock_module_0.sync_reset_por.data_sync_0_ ),
    .R(1'h1),
    .S(_00127_)
  );
  DFFSR _06504_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_reset_por.data_sync_0_ ),
    .Q( clock_module_0.por ),
    .R(1'h1),
    .S(_00128_)
  );
  INVX1 _06505_ (
    .A( dbg_0.mem_ctl_1_ ),
    .Y(_00259_)
  );
  INVX1 _06506_ (
    .A( dbg_0.mem_data_15_ ),
    .Y(_00260_)
  );
  INVX1 _06507_ (
    .A( dbg_0.mem_data_14_ ),
    .Y(_00261_)
  );
  INVX1 _06508_ (
    .A( dbg_0.mem_data_13_ ),
    .Y(_00262_)
  );
  INVX1 _06509_ (
    .A( dbg_0.mem_data_12_ ),
    .Y(_00263_)
  );
  INVX1 _06510_ (
    .A( dbg_0.mem_data_11_ ),
    .Y(_00264_)
  );
  INVX1 _06511_ (
    .A( dbg_0.mem_data_10_ ),
    .Y(_00265_)
  );
  INVX1 _06512_ (
    .A( dbg_0.mem_data_9_ ),
    .Y(_00266_)
  );
  INVX1 _06513_ (
    .A( dbg_0.mem_data_8_ ),
    .Y(_00267_)
  );
  INVX1 _06514_ (
    .A( dbg_0.mem_data_7_ ),
    .Y(_00268_)
  );
  INVX1 _06515_ (
    .A( dbg_0.mem_data_6_ ),
    .Y(_00269_)
  );
  INVX1 _06516_ (
    .A( dbg_0.mem_data_5_ ),
    .Y(_00270_)
  );
  INVX1 _06517_ (
    .A( dbg_0.mem_data_4_ ),
    .Y(_00271_)
  );
  INVX1 _06518_ (
    .A( dbg_0.mem_data_3_ ),
    .Y(_00272_)
  );
  INVX1 _06519_ (
    .A( dbg_0.mem_data_2_ ),
    .Y(_00273_)
  );
  INVX1 _06520_ (
    .A( dbg_0.mem_data_1_ ),
    .Y(_00274_)
  );
  INVX1 _06521_ (
    .A( dbg_0.mem_data_0_ ),
    .Y(_00275_)
  );
  INVX1 _06522_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00276_)
  );
  INVX1 _06523_ (
    .A( dbg_0.mem_cnt_1_ ),
    .Y(_00277_)
  );
  INVX1 _06524_ (
    .A( dbg_0.mem_cnt_0_ ),
    .Y(_00278_)
  );
  INVX1 _06525_ (
    .A( dbg_0.mem_cnt_7_ ),
    .Y(_00279_)
  );
  INVX1 _06526_ (
    .A( dbg_0.mem_start ),
    .Y(_00280_)
  );
  INVX1 _06527_ (
    .A( dbg_0.mem_startb ),
    .Y(_00281_)
  );
  INVX1 _06528_ (
    .A( dbg_0.mem_state_1_ ),
    .Y(_00282_)
  );
  INVX1 _06529_ (
    .A( dbg_0.dbg_addr_0_ ),
    .Y(_00283_)
  );
  INVX1 _06530_ (
    .A( dbg_0.dbg_mem_rd_dly ),
    .Y(_00284_)
  );
  INVX1 _06531_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00285_)
  );
  INVX1 _06532_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .Y(_00286_)
  );
  INVX1 _06533_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .Y(_00287_)
  );
  INVX1 _06534_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .Y(_00288_)
  );
  INVX1 _06535_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .Y(_00289_)
  );
  INVX1 _06536_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .Y(_00290_)
  );
  INVX1 _06537_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .Y(_00291_)
  );
  INVX1 _06538_ (
    .A( dbg_0.dbg_din_9_ ),
    .Y(_00292_)
  );
  INVX1 _06539_ (
    .A( dbg_0.dbg_din_10_ ),
    .Y(_00293_)
  );
  INVX1 _06540_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .Y(_00294_)
  );
  INVX1 _06541_ (
    .A( dbg_0.dbg_din_13_ ),
    .Y(_00295_)
  );
  INVX1 _06542_ (
    .A( dbg_0.dbg_din_15_ ),
    .Y(_00296_)
  );
  INVX1 _06543_ (
    .A(cpu_en),
    .Y(_00297_)
  );
  INVX1 _06544_ (
    .A( dbg_0.inc_step_1_ ),
    .Y(_00298_)
  );
  INVX1 _06545_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00167_)
  );
  OR2X1 _06546_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_addr_1_ ),
    .Y(_00299_)
  );
  OR2X1 _06547_ (
    .A( dbg_0.dbg_addr_0_ ),
    .B(_00299_),
    .Y(_00300_)
  );
  OR2X1 _06548_ (
    .A( dbg_0.dbg_addr_4_ ),
    .B( dbg_0.dbg_addr_5_ ),
    .Y(_00301_)
  );
  NOR2X1 _06549_ (
    .A( dbg_0.dbg_addr_3_ ),
    .B(_00301_),
    .Y(_00302_)
  );
  NAND2X1 _06550_ (
    .A( dbg_0.dbg_addr_2_ ),
    .B(_00302_),
    .Y(_00303_)
  );
  NOR2X1 _06551_ (
    .A(_00300_),
    .B(_00303_),
    .Y(_00304_)
  );
  AND2X1 _06552_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00304_),
    .Y(_00305_)
  );
  NOR2X1 _06553_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_addr_2_ ),
    .Y(_00306_)
  );
  MUX2X1 _06554_ (
    .A( dbg_0.dbg_din_3_ ),
    .B( dbg_0.dbg_i2c_0.mem_bw ),
    .S(_00305_),
    .Y(_00307_)
  );
  INVX1 _06555_ (
    .A(_00307_),
    .Y(_00258_)
  );
  MUX2X1 _06556_ (
    .A( dbg_0.dbg_din_2_ ),
    .B( dbg_0.mem_ctl_2_ ),
    .S(_00305_),
    .Y(_00308_)
  );
  INVX1 _06557_ (
    .A(_00308_),
    .Y(_00257_)
  );
  MUX2X1 _06558_ (
    .A( dbg_0.dbg_din_1_ ),
    .B( dbg_0.mem_ctl_1_ ),
    .S(_00305_),
    .Y(_00309_)
  );
  INVX1 _06559_ (
    .A(_00309_),
    .Y(_00256_)
  );
  OAI21X1 _06560_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00283_),
    .C(_00299_),
    .Y(_00310_)
  );
  AOI21X1 _06561_ (
    .A(_00276_),
    .B(_00303_),
    .C(_00310_),
    .Y(_00311_)
  );
  NAND2X1 _06562_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00311_),
    .Y(_00312_)
  );
  NAND2X1 _06563_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B( dbg_0.mem_state_1_ ),
    .Y(_00313_)
  );
  NOR2X1 _06564_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00313_),
    .Y(_00314_)
  );
  OR2X1 _06565_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00313_),
    .Y(_00315_)
  );
  OAI21X1 _06566_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00313_),
    .C(_00284_),
    .Y(_00316_)
  );
  INVX1 _06567_ (
    .A(_00316_),
    .Y(_00317_)
  );
  AOI21X1 _06568_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00311_),
    .C(_00316_),
    .Y(_00318_)
  );
  NAND2X1 _06569_ (
    .A(_00312_),
    .B(_00317_),
    .Y(_00319_)
  );
  NAND2X1 _06570_ (
    .A( dbg_0.dbg_reg_din_15_ ),
    .B(_00314_),
    .Y(_00320_)
  );
  NOR2X1 _06571_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00284_),
    .Y(_00321_)
  );
  NAND2X1 _06572_ (
    .A( dbg_0.dbg_mem_din_15_ ),
    .B(_00321_),
    .Y(_00322_)
  );
  OAI21X1 _06573_ (
    .A(_00314_),
    .B(_00322_),
    .C(_00320_),
    .Y(_00323_)
  );
  AOI22X1 _06574_ (
    .A( dbg_0.mem_data_15_ ),
    .B(_00318_),
    .C(_00323_),
    .D(_00312_),
    .Y(_00324_)
  );
  OAI21X1 _06575_ (
    .A(_00296_),
    .B(_00312_),
    .C(_00324_),
    .Y(_00255_)
  );
  NAND2X1 _06576_ (
    .A( dbg_0.dbg_reg_din_14_ ),
    .B(_00314_),
    .Y(_00325_)
  );
  NAND2X1 _06577_ (
    .A( dbg_0.dbg_mem_din_14_ ),
    .B(_00321_),
    .Y(_00326_)
  );
  OAI21X1 _06578_ (
    .A(_00314_),
    .B(_00326_),
    .C(_00325_),
    .Y(_00327_)
  );
  MUX2X1 _06579_ (
    .A(_00327_),
    .B( dbg_0.dbg_din_14_ ),
    .S(_00312_),
    .Y(_00328_)
  );
  OAI21X1 _06580_ (
    .A(_00261_),
    .B(_00319_),
    .C(_00328_),
    .Y(_00254_)
  );
  NAND2X1 _06581_ (
    .A( dbg_0.dbg_reg_din_13_ ),
    .B(_00314_),
    .Y(_00329_)
  );
  NAND2X1 _06582_ (
    .A( dbg_0.dbg_mem_din_13_ ),
    .B(_00321_),
    .Y(_00330_)
  );
  OAI21X1 _06583_ (
    .A(_00314_),
    .B(_00330_),
    .C(_00329_),
    .Y(_00331_)
  );
  AOI22X1 _06584_ (
    .A( dbg_0.mem_data_13_ ),
    .B(_00318_),
    .C(_00331_),
    .D(_00312_),
    .Y(_00332_)
  );
  OAI21X1 _06585_ (
    .A(_00295_),
    .B(_00312_),
    .C(_00332_),
    .Y(_00253_)
  );
  NAND2X1 _06586_ (
    .A( dbg_0.dbg_reg_din_12_ ),
    .B(_00314_),
    .Y(_00333_)
  );
  NAND2X1 _06587_ (
    .A( dbg_0.dbg_mem_din_12_ ),
    .B(_00321_),
    .Y(_00334_)
  );
  OAI21X1 _06588_ (
    .A(_00314_),
    .B(_00334_),
    .C(_00333_),
    .Y(_00335_)
  );
  MUX2X1 _06589_ (
    .A(_00335_),
    .B( dbg_0.dbg_din_12_ ),
    .S(_00312_),
    .Y(_00336_)
  );
  OAI21X1 _06590_ (
    .A(_00263_),
    .B(_00319_),
    .C(_00336_),
    .Y(_00252_)
  );
  NAND2X1 _06591_ (
    .A( dbg_0.dbg_reg_din_11_ ),
    .B(_00314_),
    .Y(_00337_)
  );
  NAND2X1 _06592_ (
    .A( dbg_0.dbg_mem_din_11_ ),
    .B(_00321_),
    .Y(_00338_)
  );
  OAI21X1 _06593_ (
    .A(_00314_),
    .B(_00338_),
    .C(_00337_),
    .Y(_00339_)
  );
  MUX2X1 _06594_ (
    .A(_00339_),
    .B( dbg_0.dbg_din_11_ ),
    .S(_00312_),
    .Y(_00340_)
  );
  OAI21X1 _06595_ (
    .A(_00264_),
    .B(_00319_),
    .C(_00340_),
    .Y(_00251_)
  );
  NAND2X1 _06596_ (
    .A( dbg_0.dbg_reg_din_10_ ),
    .B(_00314_),
    .Y(_00341_)
  );
  NAND2X1 _06597_ (
    .A( dbg_0.dbg_mem_din_10_ ),
    .B(_00321_),
    .Y(_00342_)
  );
  OAI21X1 _06598_ (
    .A(_00314_),
    .B(_00342_),
    .C(_00341_),
    .Y(_00343_)
  );
  AOI22X1 _06599_ (
    .A( dbg_0.mem_data_10_ ),
    .B(_00318_),
    .C(_00343_),
    .D(_00312_),
    .Y(_00344_)
  );
  OAI21X1 _06600_ (
    .A(_00293_),
    .B(_00312_),
    .C(_00344_),
    .Y(_00250_)
  );
  NAND2X1 _06601_ (
    .A( dbg_0.dbg_reg_din_9_ ),
    .B(_00314_),
    .Y(_00345_)
  );
  NAND2X1 _06602_ (
    .A( dbg_0.dbg_mem_din_9_ ),
    .B(_00321_),
    .Y(_00346_)
  );
  OAI21X1 _06603_ (
    .A(_00314_),
    .B(_00346_),
    .C(_00345_),
    .Y(_00347_)
  );
  AOI22X1 _06604_ (
    .A( dbg_0.mem_data_9_ ),
    .B(_00318_),
    .C(_00347_),
    .D(_00312_),
    .Y(_00348_)
  );
  OAI21X1 _06605_ (
    .A(_00292_),
    .B(_00312_),
    .C(_00348_),
    .Y(_00249_)
  );
  NAND2X1 _06606_ (
    .A( dbg_0.dbg_reg_din_8_ ),
    .B(_00314_),
    .Y(_00349_)
  );
  NAND2X1 _06607_ (
    .A( dbg_0.dbg_mem_din_8_ ),
    .B(_00321_),
    .Y(_00350_)
  );
  OAI21X1 _06608_ (
    .A(_00314_),
    .B(_00350_),
    .C(_00349_),
    .Y(_00351_)
  );
  MUX2X1 _06609_ (
    .A(_00351_),
    .B( dbg_0.dbg_din_8_ ),
    .S(_00312_),
    .Y(_00352_)
  );
  OAI21X1 _06610_ (
    .A(_00267_),
    .B(_00319_),
    .C(_00352_),
    .Y(_00248_)
  );
  AND2X1 _06611_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00353_)
  );
  NAND2X1 _06612_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00354_)
  );
  MUX2X1 _06613_ (
    .A( dbg_0.dbg_mem_din_7_ ),
    .B( dbg_0.dbg_mem_din_15_ ),
    .S(_00354_),
    .Y(_00355_)
  );
  AND2X1 _06614_ (
    .A(_00315_),
    .B(_00355_),
    .Y(_00356_)
  );
  OAI21X1 _06615_ (
    .A( dbg_0.dbg_reg_din_7_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00357_)
  );
  OAI21X1 _06616_ (
    .A(_00356_),
    .B(_00357_),
    .C(_00312_),
    .Y(_00358_)
  );
  OAI21X1 _06617_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00312_),
    .C(_00358_),
    .Y(_00359_)
  );
  OAI21X1 _06618_ (
    .A(_00268_),
    .B(_00319_),
    .C(_00359_),
    .Y(_00247_)
  );
  MUX2X1 _06619_ (
    .A( dbg_0.dbg_mem_din_6_ ),
    .B( dbg_0.dbg_mem_din_14_ ),
    .S(_00354_),
    .Y(_00360_)
  );
  AND2X1 _06620_ (
    .A(_00315_),
    .B(_00360_),
    .Y(_00361_)
  );
  OAI21X1 _06621_ (
    .A( dbg_0.dbg_reg_din_6_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00362_)
  );
  OAI21X1 _06622_ (
    .A(_00361_),
    .B(_00362_),
    .C(_00312_),
    .Y(_00363_)
  );
  OAI21X1 _06623_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00312_),
    .C(_00363_),
    .Y(_00364_)
  );
  OAI21X1 _06624_ (
    .A(_00269_),
    .B(_00319_),
    .C(_00364_),
    .Y(_00246_)
  );
  MUX2X1 _06625_ (
    .A( dbg_0.dbg_mem_din_5_ ),
    .B( dbg_0.dbg_mem_din_13_ ),
    .S(_00354_),
    .Y(_00365_)
  );
  AND2X1 _06626_ (
    .A(_00315_),
    .B(_00365_),
    .Y(_00366_)
  );
  OAI21X1 _06627_ (
    .A( dbg_0.dbg_reg_din_5_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00367_)
  );
  OAI21X1 _06628_ (
    .A(_00366_),
    .B(_00367_),
    .C(_00312_),
    .Y(_00368_)
  );
  OAI21X1 _06629_ (
    .A( dbg_0.dbg_din_5_ ),
    .B(_00312_),
    .C(_00368_),
    .Y(_00369_)
  );
  OAI21X1 _06630_ (
    .A(_00270_),
    .B(_00319_),
    .C(_00369_),
    .Y(_00245_)
  );
  MUX2X1 _06631_ (
    .A( dbg_0.dbg_mem_din_4_ ),
    .B( dbg_0.dbg_mem_din_12_ ),
    .S(_00354_),
    .Y(_00370_)
  );
  AND2X1 _06632_ (
    .A(_00315_),
    .B(_00370_),
    .Y(_00371_)
  );
  OAI21X1 _06633_ (
    .A( dbg_0.dbg_reg_din_4_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00372_)
  );
  OAI21X1 _06634_ (
    .A(_00371_),
    .B(_00372_),
    .C(_00312_),
    .Y(_00373_)
  );
  OAI21X1 _06635_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00312_),
    .C(_00373_),
    .Y(_00374_)
  );
  OAI21X1 _06636_ (
    .A(_00271_),
    .B(_00319_),
    .C(_00374_),
    .Y(_00244_)
  );
  MUX2X1 _06637_ (
    .A( dbg_0.dbg_mem_din_3_ ),
    .B( dbg_0.dbg_mem_din_11_ ),
    .S(_00354_),
    .Y(_00375_)
  );
  AND2X1 _06638_ (
    .A(_00315_),
    .B(_00375_),
    .Y(_00376_)
  );
  OAI21X1 _06639_ (
    .A( dbg_0.dbg_reg_din_3_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00377_)
  );
  OAI21X1 _06640_ (
    .A(_00376_),
    .B(_00377_),
    .C(_00312_),
    .Y(_00378_)
  );
  OAI21X1 _06641_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00312_),
    .C(_00378_),
    .Y(_00379_)
  );
  OAI21X1 _06642_ (
    .A(_00272_),
    .B(_00319_),
    .C(_00379_),
    .Y(_00243_)
  );
  MUX2X1 _06643_ (
    .A( dbg_0.dbg_mem_din_2_ ),
    .B( dbg_0.dbg_mem_din_10_ ),
    .S(_00354_),
    .Y(_00380_)
  );
  AND2X1 _06644_ (
    .A(_00315_),
    .B(_00380_),
    .Y(_00381_)
  );
  OAI21X1 _06645_ (
    .A( dbg_0.dbg_reg_din_2_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00382_)
  );
  OAI21X1 _06646_ (
    .A(_00381_),
    .B(_00382_),
    .C(_00312_),
    .Y(_00383_)
  );
  OAI21X1 _06647_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00312_),
    .C(_00383_),
    .Y(_00384_)
  );
  OAI21X1 _06648_ (
    .A(_00273_),
    .B(_00319_),
    .C(_00384_),
    .Y(_00242_)
  );
  MUX2X1 _06649_ (
    .A( dbg_0.dbg_mem_din_1_ ),
    .B( dbg_0.dbg_mem_din_9_ ),
    .S(_00354_),
    .Y(_00385_)
  );
  AND2X1 _06650_ (
    .A(_00315_),
    .B(_00385_),
    .Y(_00386_)
  );
  OAI21X1 _06651_ (
    .A( dbg_0.dbg_reg_din_1_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00387_)
  );
  OAI21X1 _06652_ (
    .A(_00386_),
    .B(_00387_),
    .C(_00312_),
    .Y(_00388_)
  );
  OAI21X1 _06653_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00312_),
    .C(_00388_),
    .Y(_00389_)
  );
  OAI21X1 _06654_ (
    .A(_00274_),
    .B(_00319_),
    .C(_00389_),
    .Y(_00241_)
  );
  MUX2X1 _06655_ (
    .A( dbg_0.dbg_mem_din_0_ ),
    .B( dbg_0.dbg_mem_din_8_ ),
    .S(_00354_),
    .Y(_00390_)
  );
  AND2X1 _06656_ (
    .A(_00315_),
    .B(_00390_),
    .Y(_00391_)
  );
  OAI21X1 _06657_ (
    .A( dbg_0.dbg_reg_din_0_ ),
    .B(_00315_),
    .C(_00316_),
    .Y(_00392_)
  );
  OAI21X1 _06658_ (
    .A(_00391_),
    .B(_00392_),
    .C(_00312_),
    .Y(_00393_)
  );
  OAI21X1 _06659_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00312_),
    .C(_00393_),
    .Y(_00394_)
  );
  OAI21X1 _06660_ (
    .A(_00275_),
    .B(_00319_),
    .C(_00394_),
    .Y(_00240_)
  );
  NAND2X1 _06661_ (
    .A(_00302_),
    .B(_00306_),
    .Y(_00395_)
  );
  NOR2X1 _06662_ (
    .A(_00310_),
    .B(_00395_),
    .Y(_00396_)
  );
  NAND2X1 _06663_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00396_),
    .Y(_00397_)
  );
  INVX1 _06664_ (
    .A(_00397_),
    .Y(_00398_)
  );
  OR2X1 _06665_ (
    .A( dbg_0.mem_cnt_5_ ),
    .B( dbg_0.mem_cnt_4_ ),
    .Y(_00399_)
  );
  OR2X1 _06666_ (
    .A( dbg_0.mem_cnt_7_ ),
    .B( dbg_0.mem_cnt_6_ ),
    .Y(_00400_)
  );
  NOR2X1 _06667_ (
    .A( dbg_0.mem_cnt_6_ ),
    .B(_00399_),
    .Y(_00401_)
  );
  NOR2X1 _06668_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B( dbg_0.mem_cnt_2_ ),
    .Y(_00402_)
  );
  OR2X1 _06669_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B( dbg_0.mem_cnt_3_ ),
    .Y(_00403_)
  );
  NAND2X1 _06670_ (
    .A(_00278_),
    .B(_00402_),
    .Y(_00404_)
  );
  NOR2X1 _06671_ (
    .A( dbg_0.mem_cnt_3_ ),
    .B(_00404_),
    .Y(_00405_)
  );
  NAND3X1 _06672_ (
    .A(_00279_),
    .B(_00401_),
    .C(_00405_),
    .Y(_00406_)
  );
  OR2X1 _06673_ (
    .A( dbg_0.mem_cnt_9_ ),
    .B( dbg_0.mem_cnt_8_ ),
    .Y(_00407_)
  );
  OR2X1 _06674_ (
    .A( dbg_0.mem_cnt_11_ ),
    .B( dbg_0.mem_cnt_10_ ),
    .Y(_00408_)
  );
  OR2X1 _06675_ (
    .A(_00407_),
    .B(_00408_),
    .Y(_00409_)
  );
  NOR3X1 _06676_ (
    .A( dbg_0.mem_cnt_13_ ),
    .B(_00399_),
    .C(_00400_),
    .Y(_00410_)
  );
  NOR3X1 _06677_ (
    .A( dbg_0.mem_cnt_12_ ),
    .B( dbg_0.mem_cnt_15_ ),
    .C( dbg_0.mem_cnt_14_ ),
    .Y(_00411_)
  );
  AND2X1 _06678_ (
    .A(_00402_),
    .B(_00411_),
    .Y(_00412_)
  );
  NOR3X1 _06679_ (
    .A(_00403_),
    .B(_00407_),
    .C(_00408_),
    .Y(_00413_)
  );
  NAND3X1 _06680_ (
    .A(_00410_),
    .B(_00412_),
    .C(_00413_),
    .Y(_00414_)
  );
  OAI21X1 _06681_ (
    .A(_00280_),
    .B(_00414_),
    .C(_00281_),
    .Y(_00415_)
  );
  NOR2X1 _06682_ (
    .A( dbg_0.mem_state_1_ ),
    .B( dbg_0.mem_state_0_ ),
    .Y(_00416_)
  );
  AOI22X1 _06683_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00398_),
    .C(_00415_),
    .D(_00416_),
    .Y(_00417_)
  );
  NAND2X1 _06684_ (
    .A( dbg_0.cpu_ctl_3_ ),
    .B( dbg_0.fe_mdb_in_1_ ),
    .Y(_00418_)
  );
  NOR2X1 _06685_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B( dbg_0.fe_mdb_in_5_ ),
    .Y(_00419_)
  );
  NAND3X1 _06686_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_00286_),
    .C(_00419_),
    .Y(_00420_)
  );
  NOR2X1 _06687_ (
    .A(_00418_),
    .B(_00420_),
    .Y(_00421_)
  );
  NOR2X1 _06688_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .Y(_00422_)
  );
  NAND3X1 _06689_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.decode_noirq ),
    .C(_00422_),
    .Y(_00423_)
  );
  INVX1 _06690_ (
    .A(_00423_),
    .Y(_00424_)
  );
  NOR2X1 _06691_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B( dbg_0.fe_mdb_in_13_ ),
    .Y(_00425_)
  );
  NAND3X1 _06692_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_00287_),
    .C(_00425_),
    .Y(_00426_)
  );
  NOR2X1 _06693_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_00427_)
  );
  NAND3X1 _06694_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B( dbg_0.fe_mdb_in_9_ ),
    .C(_00427_),
    .Y(_00428_)
  );
  NOR2X1 _06695_ (
    .A(_00426_),
    .B(_00428_),
    .Y(_00429_)
  );
  NAND3X1 _06696_ (
    .A(_00421_),
    .B(_00424_),
    .C(_00429_),
    .Y(_00430_)
  );
  AND2X1 _06697_ (
    .A(dbg_en),
    .B(_06327_),
    .Y(_00431_)
  );
  AOI21X1 _06698_ (
    .A( dbg_0.cpu_ctl_5_ ),
    .B(_00431_),
    .C( dbg_0.halt_flag ),
    .Y(_00432_)
  );
  NAND2X1 _06699_ (
    .A(_00430_),
    .B(_00432_),
    .Y(_00433_)
  );
  INVX1 _06700_ (
    .A(_00433_),
    .Y(_00434_)
  );
  OAI21X1 _06701_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_00417_),
    .C(_00434_),
    .Y(_00435_)
  );
  NOR2X1 _06702_ (
    .A(_00282_),
    .B( dbg_0.mem_state_0_ ),
    .Y(_00436_)
  );
  NAND2X1 _06703_ (
    .A( dbg_0.dbg_din_1_ ),
    .B( dbg_0.cpu_stat_full_0_ ),
    .Y(_00437_)
  );
  OAI21X1 _06704_ (
    .A(_00397_),
    .B(_00437_),
    .C(_00435_),
    .Y(_00438_)
  );
  NOR2X1 _06705_ (
    .A(_00436_),
    .B(_00438_),
    .Y(_00239_)
  );
  NAND2X1 _06706_ (
    .A( dbg_0.mem_start ),
    .B(_00414_),
    .Y(_00439_)
  );
  NOR2X1 _06707_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_rd_rdy ),
    .Y(_00440_)
  );
  NOR2X1 _06708_ (
    .A(_00414_),
    .B(_00440_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_end )
  );
  AOI21X1 _06709_ (
    .A(_00276_),
    .B(_00439_),
    .C( dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00238_)
  );
  MUX2X1 _06710_ (
    .A( clock_module_0.dbg_cpu_reset ),
    .B( dbg_0.dbg_din_6_ ),
    .S(_00397_),
    .Y(_00441_)
  );
  INVX1 _06711_ (
    .A(_00441_),
    .Y(_00237_)
  );
  MUX2X1 _06712_ (
    .A( dbg_0.cpu_ctl_5_ ),
    .B( dbg_0.dbg_din_5_ ),
    .S(_00397_),
    .Y(_00442_)
  );
  INVX1 _06713_ (
    .A(_00442_),
    .Y(_00236_)
  );
  MUX2X1 _06714_ (
    .A( dbg_0.cpu_ctl_4_ ),
    .B( dbg_0.dbg_din_4_ ),
    .S(_00397_),
    .Y(_00443_)
  );
  INVX1 _06715_ (
    .A(_00443_),
    .Y(_00235_)
  );
  MUX2X1 _06716_ (
    .A( dbg_0.cpu_ctl_3_ ),
    .B( dbg_0.dbg_din_3_ ),
    .S(_00397_),
    .Y(_00444_)
  );
  INVX1 _06717_ (
    .A(_00444_),
    .Y(_00234_)
  );
  AOI21X1 _06718_ (
    .A( dbg_0.mem_state_0_ ),
    .B( dbg_0.cpu_stat_full_0_ ),
    .C( dbg_0.mem_state_1_ ),
    .Y(_00445_)
  );
  OAI21X1 _06719_ (
    .A( dbg_0.mem_state_0_ ),
    .B(_00415_),
    .C(_00445_),
    .Y(_00446_)
  );
  INVX1 _06720_ (
    .A(_00446_),
    .Y( dbg_0.mem_state_nxt_0_ )
  );
  NOR2X1 _06721_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B(_00282_),
    .Y( dbg_0.dbg_mem_en )
  );
  AND2X1 _06722_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B( dbg_0.mem_state_1_ ),
    .Y(_00447_)
  );
  NAND2X1 _06723_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B( dbg_0.dbg_mem_en ),
    .Y(_00448_)
  );
  NOR2X1 _06724_ (
    .A(_00353_),
    .B(_00448_),
    .Y( dbg_0.dbg_mem_wr_0_ )
  );
  AOI21X1 _06725_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00285_),
    .C(_00448_),
    .Y( dbg_0.dbg_mem_wr_1_ )
  );
  OAI21X1 _06726_ (
    .A( dbg_0.mem_state_0_ ),
    .B(_00415_),
    .C( dbg_0.cpu_stat_full_0_ ),
    .Y(_00449_)
  );
  NOR2X1 _06727_ (
    .A( dbg_0.mem_state_1_ ),
    .B(_00449_),
    .Y( dbg_0.mem_state_nxt_1_ )
  );
  NOR2X1 _06728_ (
    .A(_00259_),
    .B(_00313_),
    .Y( dbg_0.dbg_reg_wr )
  );
  OR2X1 _06729_ (
    .A(_00283_),
    .B(_00299_),
    .Y(_00450_)
  );
  NOR2X1 _06730_ (
    .A(_00303_),
    .B(_00450_),
    .Y(_00451_)
  );
  AND2X1 _06731_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00451_),
    .Y(_00452_)
  );
  NAND2X1 _06732_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00451_),
    .Y(_00453_)
  );
  NOR2X1 _06733_ (
    .A( dbg_0.dbg_rd_rdy ),
    .B(_00447_),
    .Y(_00454_)
  );
  NOR2X1 _06734_ (
    .A(_00276_),
    .B(_00454_),
    .Y(_00455_)
  );
  OAI21X1 _06735_ (
    .A( dbg_0.dbg_rd_rdy ),
    .B(_00447_),
    .C( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00456_)
  );
  AND2X1 _06736_ (
    .A(_00414_),
    .B(_00455_),
    .Y(_00457_)
  );
  NAND2X1 _06737_ (
    .A(_00414_),
    .B(_00455_),
    .Y(_00458_)
  );
  OR2X1 _06738_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.mem_ctl_2_ ),
    .Y(_00459_)
  );
  NOR2X1 _06739_ (
    .A(_00456_),
    .B(_00459_),
    .Y(_00460_)
  );
  NAND3X1 _06740_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .B(_00457_),
    .C(_00459_),
    .Y(_00461_)
  );
  OAI21X1 _06741_ (
    .A(_00458_),
    .B(_00460_),
    .C(_00285_),
    .Y(_00462_)
  );
  NAND2X1 _06742_ (
    .A(_00461_),
    .B(_00462_),
    .Y(_00463_)
  );
  NAND2X1 _06743_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00452_),
    .Y(_00464_)
  );
  OAI21X1 _06744_ (
    .A(_00452_),
    .B(_00463_),
    .C(_00464_),
    .Y(_00133_)
  );
  AND2X1 _06745_ (
    .A(_00414_),
    .B(_00460_),
    .Y(_00465_)
  );
  NAND2X1 _06746_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .B(_00465_),
    .Y(_00466_)
  );
  XNOR2X1 _06747_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .B(_00465_),
    .Y(_00467_)
  );
  XNOR2X1 _06748_ (
    .A(_00461_),
    .B(_00467_),
    .Y(_00468_)
  );
  NAND2X1 _06749_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00452_),
    .Y(_00469_)
  );
  OAI21X1 _06750_ (
    .A(_00452_),
    .B(_00468_),
    .C(_00469_),
    .Y(_00140_)
  );
  OAI21X1 _06751_ (
    .A(_00461_),
    .B(_00467_),
    .C(_00466_),
    .Y(_00470_)
  );
  AND2X1 _06752_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00470_),
    .Y(_00471_)
  );
  NAND2X1 _06753_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00470_),
    .Y(_00472_)
  );
  OAI21X1 _06754_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00470_),
    .C(_00453_),
    .Y(_00473_)
  );
  NAND2X1 _06755_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00452_),
    .Y(_00474_)
  );
  OAI21X1 _06756_ (
    .A(_00471_),
    .B(_00473_),
    .C(_00474_),
    .Y(_00141_)
  );
  NAND3X1 _06757_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_3_ ),
    .C(_00470_),
    .Y(_00475_)
  );
  XOR2X1 _06758_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_00472_),
    .Y(_00476_)
  );
  NAND2X1 _06759_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00452_),
    .Y(_00477_)
  );
  OAI21X1 _06760_ (
    .A(_00452_),
    .B(_00476_),
    .C(_00477_),
    .Y(_00142_)
  );
  NOR2X1 _06761_ (
    .A(_00288_),
    .B(_00475_),
    .Y(_00478_)
  );
  XNOR2X1 _06762_ (
    .A(_00288_),
    .B(_00475_),
    .Y(_00479_)
  );
  NAND2X1 _06763_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00452_),
    .Y(_00480_)
  );
  OAI21X1 _06764_ (
    .A(_00452_),
    .B(_00479_),
    .C(_00480_),
    .Y(_00143_)
  );
  NAND2X1 _06765_ (
    .A( dbg_0.dbg_din_5_ ),
    .B(_00452_),
    .Y(_00481_)
  );
  NOR3X1 _06766_ (
    .A(_00288_),
    .B(_00289_),
    .C(_00475_),
    .Y(_00482_)
  );
  XNOR2X1 _06767_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .B(_00478_),
    .Y(_00483_)
  );
  OAI21X1 _06768_ (
    .A(_00452_),
    .B(_00483_),
    .C(_00481_),
    .Y(_00144_)
  );
  NAND2X1 _06769_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00452_),
    .Y(_00484_)
  );
  AND2X1 _06770_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00482_),
    .Y(_00485_)
  );
  OAI21X1 _06771_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00482_),
    .C(_00453_),
    .Y(_00486_)
  );
  OAI21X1 _06772_ (
    .A(_00485_),
    .B(_00486_),
    .C(_00484_),
    .Y(_00145_)
  );
  NAND2X1 _06773_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00452_),
    .Y(_00487_)
  );
  NAND3X1 _06774_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B( dbg_0.dbg_mem_addr_7_ ),
    .C(_00482_),
    .Y(_00488_)
  );
  INVX1 _06775_ (
    .A(_00488_),
    .Y(_00489_)
  );
  OAI21X1 _06776_ (
    .A( dbg_0.dbg_mem_addr_7_ ),
    .B(_00485_),
    .C(_00453_),
    .Y(_00490_)
  );
  OAI21X1 _06777_ (
    .A(_00489_),
    .B(_00490_),
    .C(_00487_),
    .Y(_00146_)
  );
  NAND2X1 _06778_ (
    .A( dbg_0.dbg_din_8_ ),
    .B(_00452_),
    .Y(_00491_)
  );
  XNOR2X1 _06779_ (
    .A(_00290_),
    .B(_00488_),
    .Y(_00492_)
  );
  OAI21X1 _06780_ (
    .A(_00452_),
    .B(_00492_),
    .C(_00491_),
    .Y(_00147_)
  );
  OAI21X1 _06781_ (
    .A(_00290_),
    .B(_00488_),
    .C(_00291_),
    .Y(_00493_)
  );
  NOR3X1 _06782_ (
    .A(_00290_),
    .B(_00291_),
    .C(_00488_),
    .Y(_00494_)
  );
  NOR2X1 _06783_ (
    .A(_00452_),
    .B(_00494_),
    .Y(_00495_)
  );
  NAND2X1 _06784_ (
    .A(_00493_),
    .B(_00495_),
    .Y(_00496_)
  );
  OAI21X1 _06785_ (
    .A(_00292_),
    .B(_00453_),
    .C(_00496_),
    .Y(_00148_)
  );
  NAND2X1 _06786_ (
    .A( dbg_0.dbg_din_10_ ),
    .B(_00452_),
    .Y(_00497_)
  );
  NAND2X1 _06787_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00494_),
    .Y(_00498_)
  );
  XNOR2X1 _06788_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00494_),
    .Y(_00499_)
  );
  OAI21X1 _06789_ (
    .A(_00452_),
    .B(_00499_),
    .C(_00497_),
    .Y(_00134_)
  );
  NAND2X1 _06790_ (
    .A( dbg_0.dbg_din_11_ ),
    .B(_00452_),
    .Y(_00500_)
  );
  NAND3X1 _06791_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B( dbg_0.dbg_mem_addr_11_ ),
    .C(_00494_),
    .Y(_00501_)
  );
  XOR2X1 _06792_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .B(_00498_),
    .Y(_00502_)
  );
  OAI21X1 _06793_ (
    .A(_00452_),
    .B(_00502_),
    .C(_00500_),
    .Y(_00135_)
  );
  NAND2X1 _06794_ (
    .A( dbg_0.dbg_din_12_ ),
    .B(_00452_),
    .Y(_00503_)
  );
  NOR2X1 _06795_ (
    .A(_00294_),
    .B(_00501_),
    .Y(_00504_)
  );
  XNOR2X1 _06796_ (
    .A(_00294_),
    .B(_00501_),
    .Y(_00505_)
  );
  OAI21X1 _06797_ (
    .A(_00452_),
    .B(_00505_),
    .C(_00503_),
    .Y(_00136_)
  );
  NAND2X1 _06798_ (
    .A( dbg_0.dbg_din_13_ ),
    .B(_00452_),
    .Y(_00506_)
  );
  NAND2X1 _06799_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00504_),
    .Y(_00507_)
  );
  XNOR2X1 _06800_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00504_),
    .Y(_00508_)
  );
  OAI21X1 _06801_ (
    .A(_00452_),
    .B(_00508_),
    .C(_00506_),
    .Y(_00137_)
  );
  NAND2X1 _06802_ (
    .A( dbg_0.dbg_din_14_ ),
    .B(_00452_),
    .Y(_00509_)
  );
  NAND3X1 _06803_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B( dbg_0.dbg_mem_addr_14_ ),
    .C(_00504_),
    .Y(_00510_)
  );
  XOR2X1 _06804_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_00507_),
    .Y(_00511_)
  );
  OAI21X1 _06805_ (
    .A(_00452_),
    .B(_00511_),
    .C(_00509_),
    .Y(_00138_)
  );
  XOR2X1 _06806_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B(_00510_),
    .Y(_00512_)
  );
  MUX2X1 _06807_ (
    .A(_00296_),
    .B(_00512_),
    .S(_00452_),
    .Y(_00139_)
  );
  NAND3X1 _06808_ (
    .A(_00276_),
    .B( dbg_0.dbg_addr_0_ ),
    .C( dbg_0.dbg_addr_1_ ),
    .Y(_00513_)
  );
  NOR2X1 _06809_ (
    .A(_00303_),
    .B(_00513_),
    .Y(_00514_)
  );
  AND2X1 _06810_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00514_),
    .Y(_00515_)
  );
  NAND2X1 _06811_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00514_),
    .Y(_00516_)
  );
  XNOR2X1 _06812_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B(_00457_),
    .Y(_00517_)
  );
  NAND2X1 _06813_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00515_),
    .Y(_00518_)
  );
  OAI21X1 _06814_ (
    .A(_00515_),
    .B(_00517_),
    .C(_00518_),
    .Y(_00149_)
  );
  NAND3X1 _06815_ (
    .A(_00277_),
    .B(_00278_),
    .C(_00457_),
    .Y(_00519_)
  );
  OAI21X1 _06816_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B(_00458_),
    .C( dbg_0.mem_cnt_1_ ),
    .Y(_00520_)
  );
  AND2X1 _06817_ (
    .A(_00519_),
    .B(_00520_),
    .Y(_00521_)
  );
  NAND2X1 _06818_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00515_),
    .Y(_00522_)
  );
  OAI21X1 _06819_ (
    .A(_00515_),
    .B(_00521_),
    .C(_00522_),
    .Y(_00156_)
  );
  XOR2X1 _06820_ (
    .A( dbg_0.mem_cnt_2_ ),
    .B(_00519_),
    .Y(_00523_)
  );
  NAND2X1 _06821_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00515_),
    .Y(_00524_)
  );
  OAI21X1 _06822_ (
    .A(_00515_),
    .B(_00523_),
    .C(_00524_),
    .Y(_00157_)
  );
  OAI21X1 _06823_ (
    .A(_00404_),
    .B(_00458_),
    .C( dbg_0.mem_cnt_3_ ),
    .Y(_00525_)
  );
  NAND2X1 _06824_ (
    .A(_00405_),
    .B(_00457_),
    .Y(_00526_)
  );
  NAND3X1 _06825_ (
    .A(_00516_),
    .B(_00525_),
    .C(_00526_),
    .Y(_00527_)
  );
  OAI21X1 _06826_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00516_),
    .C(_00527_),
    .Y(_00528_)
  );
  INVX1 _06827_ (
    .A(_00528_),
    .Y(_00158_)
  );
  XOR2X1 _06828_ (
    .A( dbg_0.mem_cnt_4_ ),
    .B(_00526_),
    .Y(_00529_)
  );
  NAND2X1 _06829_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00515_),
    .Y(_00530_)
  );
  OAI21X1 _06830_ (
    .A(_00515_),
    .B(_00529_),
    .C(_00530_),
    .Y(_00159_)
  );
  OR2X1 _06831_ (
    .A(_00399_),
    .B(_00526_),
    .Y(_00531_)
  );
  OAI21X1 _06832_ (
    .A( dbg_0.mem_cnt_4_ ),
    .B(_00526_),
    .C( dbg_0.mem_cnt_5_ ),
    .Y(_00532_)
  );
  AND2X1 _06833_ (
    .A(_00531_),
    .B(_00532_),
    .Y(_00533_)
  );
  NAND2X1 _06834_ (
    .A( dbg_0.dbg_din_5_ ),
    .B(_00515_),
    .Y(_00534_)
  );
  OAI21X1 _06835_ (
    .A(_00515_),
    .B(_00533_),
    .C(_00534_),
    .Y(_00160_)
  );
  XOR2X1 _06836_ (
    .A( dbg_0.mem_cnt_6_ ),
    .B(_00531_),
    .Y(_00535_)
  );
  NOR2X1 _06837_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00516_),
    .Y(_00536_)
  );
  AOI21X1 _06838_ (
    .A(_00516_),
    .B(_00535_),
    .C(_00536_),
    .Y(_00161_)
  );
  OAI21X1 _06839_ (
    .A( dbg_0.mem_cnt_6_ ),
    .B(_00531_),
    .C( dbg_0.mem_cnt_7_ ),
    .Y(_00537_)
  );
  OR2X1 _06840_ (
    .A(_00406_),
    .B(_00458_),
    .Y(_00538_)
  );
  AND2X1 _06841_ (
    .A(_00537_),
    .B(_00538_),
    .Y(_00539_)
  );
  NAND2X1 _06842_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00515_),
    .Y(_00540_)
  );
  OAI21X1 _06843_ (
    .A(_00515_),
    .B(_00539_),
    .C(_00540_),
    .Y(_00162_)
  );
  XOR2X1 _06844_ (
    .A( dbg_0.mem_cnt_8_ ),
    .B(_00538_),
    .Y(_00541_)
  );
  NAND2X1 _06845_ (
    .A( dbg_0.dbg_din_8_ ),
    .B(_00515_),
    .Y(_00542_)
  );
  OAI21X1 _06846_ (
    .A(_00515_),
    .B(_00541_),
    .C(_00542_),
    .Y(_00163_)
  );
  OR2X1 _06847_ (
    .A(_00407_),
    .B(_00538_),
    .Y(_00543_)
  );
  OAI21X1 _06848_ (
    .A( dbg_0.mem_cnt_8_ ),
    .B(_00538_),
    .C( dbg_0.mem_cnt_9_ ),
    .Y(_00544_)
  );
  AND2X1 _06849_ (
    .A(_00543_),
    .B(_00544_),
    .Y(_00545_)
  );
  NAND2X1 _06850_ (
    .A( dbg_0.dbg_din_9_ ),
    .B(_00515_),
    .Y(_00546_)
  );
  OAI21X1 _06851_ (
    .A(_00515_),
    .B(_00545_),
    .C(_00546_),
    .Y(_00164_)
  );
  OAI21X1 _06852_ (
    .A(_00407_),
    .B(_00538_),
    .C( dbg_0.mem_cnt_10_ ),
    .Y(_00547_)
  );
  NOR2X1 _06853_ (
    .A( dbg_0.mem_cnt_10_ ),
    .B(_00543_),
    .Y(_00548_)
  );
  NOR2X1 _06854_ (
    .A(_00515_),
    .B(_00548_),
    .Y(_00549_)
  );
  AOI22X1 _06855_ (
    .A(_00293_),
    .B(_00515_),
    .C(_00547_),
    .D(_00549_),
    .Y(_00150_)
  );
  XNOR2X1 _06856_ (
    .A( dbg_0.mem_cnt_11_ ),
    .B(_00548_),
    .Y(_00550_)
  );
  NAND2X1 _06857_ (
    .A( dbg_0.dbg_din_11_ ),
    .B(_00515_),
    .Y(_00551_)
  );
  OAI21X1 _06858_ (
    .A(_00515_),
    .B(_00550_),
    .C(_00551_),
    .Y(_00151_)
  );
  NAND2X1 _06859_ (
    .A( dbg_0.mem_cnt_12_ ),
    .B(_00455_),
    .Y(_00552_)
  );
  XNOR2X1 _06860_ (
    .A( dbg_0.mem_cnt_12_ ),
    .B(_00457_),
    .Y(_00553_)
  );
  OAI21X1 _06861_ (
    .A(_00406_),
    .B(_00409_),
    .C(_00455_),
    .Y(_00554_)
  );
  XNOR2X1 _06862_ (
    .A(_00553_),
    .B(_00554_),
    .Y(_00555_)
  );
  NAND2X1 _06863_ (
    .A( dbg_0.dbg_din_12_ ),
    .B(_00515_),
    .Y(_00556_)
  );
  OAI21X1 _06864_ (
    .A(_00515_),
    .B(_00555_),
    .C(_00556_),
    .Y(_00152_)
  );
  OAI21X1 _06865_ (
    .A(_00553_),
    .B(_00554_),
    .C(_00552_),
    .Y(_00557_)
  );
  XNOR2X1 _06866_ (
    .A( dbg_0.mem_cnt_13_ ),
    .B(_00458_),
    .Y(_00558_)
  );
  XNOR2X1 _06867_ (
    .A(_00557_),
    .B(_00558_),
    .Y(_00559_)
  );
  MUX2X1 _06868_ (
    .A(_00295_),
    .B(_00559_),
    .S(_00515_),
    .Y(_00153_)
  );
  NAND2X1 _06869_ (
    .A( dbg_0.mem_cnt_14_ ),
    .B(_00455_),
    .Y(_00560_)
  );
  XNOR2X1 _06870_ (
    .A( dbg_0.mem_cnt_14_ ),
    .B(_00457_),
    .Y(_00561_)
  );
  AOI21X1 _06871_ (
    .A( dbg_0.mem_cnt_13_ ),
    .B(_00457_),
    .C(_00557_),
    .Y(_00562_)
  );
  XNOR2X1 _06872_ (
    .A(_00561_),
    .B(_00562_),
    .Y(_00563_)
  );
  NAND2X1 _06873_ (
    .A( dbg_0.dbg_din_14_ ),
    .B(_00515_),
    .Y(_00564_)
  );
  OAI21X1 _06874_ (
    .A(_00515_),
    .B(_00563_),
    .C(_00564_),
    .Y(_00154_)
  );
  OAI21X1 _06875_ (
    .A(_00561_),
    .B(_00562_),
    .C(_00560_),
    .Y(_00565_)
  );
  XNOR2X1 _06876_ (
    .A( dbg_0.mem_cnt_15_ ),
    .B(_00458_),
    .Y(_00566_)
  );
  OR2X1 _06877_ (
    .A(_00565_),
    .B(_00566_),
    .Y(_00567_)
  );
  OAI21X1 _06878_ (
    .A( dbg_0.mem_cnt_15_ ),
    .B(_00458_),
    .C(_00567_),
    .Y(_00568_)
  );
  NAND2X1 _06879_ (
    .A( dbg_0.dbg_din_15_ ),
    .B(_00515_),
    .Y(_00569_)
  );
  OAI21X1 _06880_ (
    .A(_00515_),
    .B(_00568_),
    .C(_00569_),
    .Y(_00155_)
  );
  NOR2X1 _06881_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00439_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_rd )
  );
  OAI21X1 _06882_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00439_),
    .C(_00276_),
    .Y(_00570_)
  );
  OAI21X1 _06883_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_i2c_0.mem_burst_rd ),
    .C(_00317_),
    .Y(_00571_)
  );
  OAI21X1 _06884_ (
    .A( dbg_0.dbg_i2c_0.dbg_rd ),
    .B(_00570_),
    .C(_00571_),
    .Y(_00572_)
  );
  INVX1 _06885_ (
    .A(_00572_),
    .Y(_00131_)
  );
  NAND2X1 _06886_ (
    .A( dbg_0.dbg_din_2_ ),
    .B( dbg_0.cpu_stat_full_0_ ),
    .Y(_00573_)
  );
  NOR2X1 _06887_ (
    .A(_00397_),
    .B(_00573_),
    .Y( dbg_0.istep )
  );
  OR2X1 _06888_ (
    .A( dbg_0.inc_step_0_ ),
    .B( dbg_0.istep ),
    .Y(_00132_)
  );
  NOR2X1 _06889_ (
    .A(_00275_),
    .B(_00353_),
    .Y(_06309_)
  );
  NOR2X1 _06890_ (
    .A(_00274_),
    .B(_00353_),
    .Y(_06316_)
  );
  NOR2X1 _06891_ (
    .A(_00273_),
    .B(_00353_),
    .Y(_06317_)
  );
  NOR2X1 _06892_ (
    .A(_00272_),
    .B(_00353_),
    .Y(_06318_)
  );
  NOR2X1 _06893_ (
    .A(_00271_),
    .B(_00353_),
    .Y(_06319_)
  );
  NOR2X1 _06894_ (
    .A(_00270_),
    .B(_00353_),
    .Y(_06320_)
  );
  NOR2X1 _06895_ (
    .A(_00269_),
    .B(_00353_),
    .Y(_06321_)
  );
  NOR2X1 _06896_ (
    .A(_00268_),
    .B(_00353_),
    .Y(_06322_)
  );
  OAI22X1 _06897_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00267_),
    .C(_00275_),
    .D(_00354_),
    .Y(_06323_)
  );
  OAI22X1 _06898_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00266_),
    .C(_00274_),
    .D(_00354_),
    .Y(_06324_)
  );
  OAI22X1 _06899_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00265_),
    .C(_00273_),
    .D(_00354_),
    .Y(_06310_)
  );
  OAI22X1 _06900_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00264_),
    .C(_00272_),
    .D(_00354_),
    .Y(_06311_)
  );
  OAI22X1 _06901_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00263_),
    .C(_00271_),
    .D(_00354_),
    .Y(_06312_)
  );
  OAI22X1 _06902_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00262_),
    .C(_00270_),
    .D(_00354_),
    .Y(_06313_)
  );
  OAI22X1 _06903_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00261_),
    .C(_00269_),
    .D(_00354_),
    .Y(_06314_)
  );
  OAI22X1 _06904_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00260_),
    .C(_00268_),
    .D(_00354_),
    .Y(_06315_)
  );
  NOR2X1 _06905_ (
    .A(_00395_),
    .B(_00513_),
    .Y(_00574_)
  );
  NAND3X1 _06906_ (
    .A( dbg_0.dbg_din_2_ ),
    .B( dbg_0.dbg_i2c_0.dbg_wr ),
    .C(_00574_),
    .Y(_00575_)
  );
  AOI21X1 _06907_ (
    .A( dbg_0.cpu_stat_2_ ),
    .B(_00575_),
    .C(_06327_),
    .Y(_00576_)
  );
  INVX1 _06908_ (
    .A(_00576_),
    .Y(_00129_)
  );
  NAND3X1 _06909_ (
    .A( dbg_0.dbg_din_3_ ),
    .B( dbg_0.dbg_i2c_0.dbg_wr ),
    .C(_00574_),
    .Y(_00577_)
  );
  NAND2X1 _06910_ (
    .A( dbg_0.cpu_stat_3_ ),
    .B(_00577_),
    .Y(_00578_)
  );
  NAND2X1 _06911_ (
    .A(_00430_),
    .B(_00578_),
    .Y(_00130_)
  );
  AND2X1 _06912_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00305_),
    .Y(_00165_)
  );
  NAND2X1 _06913_ (
    .A( dbg_0.dbg_addr_3_ ),
    .B( dbg_0.dbg_addr_4_ ),
    .Y(_00579_)
  );
  NOR2X1 _06914_ (
    .A( dbg_0.dbg_addr_5_ ),
    .B(_00579_),
    .Y(_00580_)
  );
  NAND2X1 _06915_ (
    .A(_00306_),
    .B(_00580_),
    .Y(_00581_)
  );
  NOR2X1 _06916_ (
    .A(_00300_),
    .B(_00581_),
    .Y(_00582_)
  );
  NOR2X1 _06917_ (
    .A(_00395_),
    .B(_00450_),
    .Y(_00583_)
  );
  NOR2X1 _06918_ (
    .A(_00300_),
    .B(_00395_),
    .Y(_00584_)
  );
  AOI22X1 _06919_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .B(_00451_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_0_ ),
    .Y(_00585_)
  );
  INVX1 _06920_ (
    .A(_00585_),
    .Y(_00586_)
  );
  AOI21X1 _06921_ (
    .A( dbg_0.mem_data_0_ ),
    .B(_00311_),
    .C(_00586_),
    .Y(_00587_)
  );
  AOI22X1 _06922_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h1),
    .Y(_00588_)
  );
  AOI22X1 _06923_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_00574_),
    .C(_00583_),
    .D(1'h1),
    .Y(_00589_)
  );
  NAND3X1 _06924_ (
    .A(_00587_),
    .B(_00588_),
    .C(_00589_),
    .Y( dbg_0.dbg_dout_0_ )
  );
  AOI22X1 _06925_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00590_)
  );
  AOI22X1 _06926_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B(_00514_),
    .C(_00584_),
    .D(1'h1),
    .Y(_00591_)
  );
  AOI22X1 _06927_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00304_),
    .C(_00451_),
    .D( dbg_0.dbg_mem_addr_1_ ),
    .Y(_00592_)
  );
  INVX1 _06928_ (
    .A(_00592_),
    .Y(_00593_)
  );
  AOI21X1 _06929_ (
    .A( dbg_0.mem_data_1_ ),
    .B(_00311_),
    .C(_00593_),
    .Y(_00594_)
  );
  NAND3X1 _06930_ (
    .A(_00590_),
    .B(_00591_),
    .C(_00594_),
    .Y( dbg_0.dbg_dout_1_ )
  );
  NAND2X1 _06931_ (
    .A( dbg_0.cpu_stat_2_ ),
    .B(_00574_),
    .Y(_00595_)
  );
  AOI22X1 _06932_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00596_)
  );
  AOI22X1 _06933_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B(_00304_),
    .C(_00451_),
    .D( dbg_0.dbg_mem_addr_2_ ),
    .Y(_00597_)
  );
  AOI22X1 _06934_ (
    .A( dbg_0.mem_cnt_2_ ),
    .B(_00514_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00598_)
  );
  NAND2X1 _06935_ (
    .A(_00597_),
    .B(_00598_),
    .Y(_00599_)
  );
  AOI21X1 _06936_ (
    .A( dbg_0.mem_data_2_ ),
    .B(_00311_),
    .C(_00599_),
    .Y(_00600_)
  );
  NAND3X1 _06937_ (
    .A(_00595_),
    .B(_00596_),
    .C(_00600_),
    .Y( dbg_0.dbg_dout_2_ )
  );
  AOI22X1 _06938_ (
    .A(1'h0),
    .B(_00583_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00601_)
  );
  AOI22X1 _06939_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00304_),
    .C(_00396_),
    .D( dbg_0.cpu_ctl_3_ ),
    .Y(_00602_)
  );
  AOI22X1 _06940_ (
    .A( dbg_0.cpu_stat_3_ ),
    .B(_00574_),
    .C(_00582_),
    .D(1'h0),
    .Y(_00603_)
  );
  AOI22X1 _06941_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_00451_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_3_ ),
    .Y(_00604_)
  );
  NAND2X1 _06942_ (
    .A(_00603_),
    .B(_00604_),
    .Y(_00605_)
  );
  AOI21X1 _06943_ (
    .A( dbg_0.mem_data_3_ ),
    .B(_00311_),
    .C(_00605_),
    .Y(_00606_)
  );
  NAND3X1 _06944_ (
    .A(_00601_),
    .B(_00602_),
    .C(_00606_),
    .Y( dbg_0.dbg_dout_3_ )
  );
  AOI22X1 _06945_ (
    .A( dbg_0.cpu_ctl_4_ ),
    .B(_00396_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00607_)
  );
  AOI22X1 _06946_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .B(_00451_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_4_ ),
    .Y(_00608_)
  );
  INVX1 _06947_ (
    .A(_00608_),
    .Y(_00609_)
  );
  AOI21X1 _06948_ (
    .A( dbg_0.mem_data_4_ ),
    .B(_00311_),
    .C(_00609_),
    .Y(_00610_)
  );
  AOI22X1 _06949_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00611_)
  );
  NAND3X1 _06950_ (
    .A(_00607_),
    .B(_00610_),
    .C(_00611_),
    .Y( dbg_0.dbg_dout_4_ )
  );
  AOI22X1 _06951_ (
    .A( dbg_0.cpu_ctl_5_ ),
    .B(_00396_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_5_ ),
    .Y(_00612_)
  );
  AOI22X1 _06952_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00613_)
  );
  AOI22X1 _06953_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00614_)
  );
  INVX1 _06954_ (
    .A(_00614_),
    .Y(_00615_)
  );
  AOI21X1 _06955_ (
    .A( dbg_0.mem_data_5_ ),
    .B(_00311_),
    .C(_00615_),
    .Y(_00616_)
  );
  NAND3X1 _06956_ (
    .A(_00612_),
    .B(_00613_),
    .C(_00616_),
    .Y( dbg_0.dbg_dout_5_ )
  );
  AOI22X1 _06957_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00451_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_6_ ),
    .Y(_00617_)
  );
  INVX1 _06958_ (
    .A(_00617_),
    .Y(_00618_)
  );
  AOI21X1 _06959_ (
    .A( dbg_0.mem_data_6_ ),
    .B(_00311_),
    .C(_00618_),
    .Y(_00619_)
  );
  AOI22X1 _06960_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00620_)
  );
  AOI22X1 _06961_ (
    .A( clock_module_0.dbg_cpu_reset ),
    .B(_00396_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00621_)
  );
  NAND3X1 _06962_ (
    .A(_00619_),
    .B(_00620_),
    .C(_00621_),
    .Y( dbg_0.dbg_dout_6_ )
  );
  AOI22X1 _06963_ (
    .A( dbg_0.mem_data_7_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_7_ ),
    .Y(_00622_)
  );
  AOI22X1 _06964_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00623_)
  );
  AOI22X1 _06965_ (
    .A( dbg_0.dbg_mem_addr_7_ ),
    .B(_00451_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00624_)
  );
  NAND3X1 _06966_ (
    .A(_00622_),
    .B(_00623_),
    .C(_00624_),
    .Y( dbg_0.dbg_dout_7_ )
  );
  AOI22X1 _06967_ (
    .A( dbg_0.mem_data_8_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_8_ ),
    .Y(_00625_)
  );
  AOI22X1 _06968_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h1),
    .Y(_00626_)
  );
  AOI22X1 _06969_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00627_)
  );
  NAND3X1 _06970_ (
    .A(_00625_),
    .B(_00626_),
    .C(_00627_),
    .Y( dbg_0.dbg_dout_8_ )
  );
  AOI22X1 _06971_ (
    .A( dbg_0.mem_data_9_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_9_ ),
    .Y(_00628_)
  );
  AOI22X1 _06972_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00629_)
  );
  AOI22X1 _06973_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .B(_00451_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00630_)
  );
  NAND3X1 _06974_ (
    .A(_00628_),
    .B(_00629_),
    .C(_00630_),
    .Y( dbg_0.dbg_dout_9_ )
  );
  AOI22X1 _06975_ (
    .A( dbg_0.mem_data_10_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_10_ ),
    .Y(_00631_)
  );
  AOI22X1 _06976_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00632_)
  );
  AOI22X1 _06977_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00451_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00633_)
  );
  NAND3X1 _06978_ (
    .A(_00631_),
    .B(_00632_),
    .C(_00633_),
    .Y( dbg_0.dbg_dout_10_ )
  );
  NAND2X1 _06979_ (
    .A(1'h0),
    .B(_00583_),
    .Y(_00634_)
  );
  AOI22X1 _06980_ (
    .A( dbg_0.mem_data_11_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_11_ ),
    .Y(_00635_)
  );
  AOI22X1 _06981_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00636_)
  );
  NAND2X1 _06982_ (
    .A(_00634_),
    .B(_00636_),
    .Y(_00637_)
  );
  AOI21X1 _06983_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .B(_00451_),
    .C(_00637_),
    .Y(_00638_)
  );
  NAND2X1 _06984_ (
    .A(_00635_),
    .B(_00638_),
    .Y( dbg_0.dbg_dout_11_ )
  );
  AOI22X1 _06985_ (
    .A( dbg_0.mem_data_12_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_12_ ),
    .Y(_00639_)
  );
  AOI22X1 _06986_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00640_)
  );
  AOI22X1 _06987_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00641_)
  );
  NAND3X1 _06988_ (
    .A(_00639_),
    .B(_00640_),
    .C(_00641_),
    .Y( dbg_0.dbg_dout_12_ )
  );
  AOI22X1 _06989_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00642_)
  );
  INVX1 _06990_ (
    .A(_00642_),
    .Y(_00643_)
  );
  AOI21X1 _06991_ (
    .A( dbg_0.mem_cnt_13_ ),
    .B(_00514_),
    .C(_00643_),
    .Y(_00644_)
  );
  AOI22X1 _06992_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00645_)
  );
  NAND2X1 _06993_ (
    .A( dbg_0.mem_data_13_ ),
    .B(_00311_),
    .Y(_00646_)
  );
  NAND3X1 _06994_ (
    .A(_00644_),
    .B(_00645_),
    .C(_00646_),
    .Y( dbg_0.dbg_dout_13_ )
  );
  AOI22X1 _06995_ (
    .A( dbg_0.mem_data_14_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_14_ ),
    .Y(_00647_)
  );
  AOI22X1 _06996_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h0),
    .Y(_00648_)
  );
  AOI22X1 _06997_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h1),
    .Y(_00649_)
  );
  NAND3X1 _06998_ (
    .A(_00647_),
    .B(_00648_),
    .C(_00649_),
    .Y( dbg_0.dbg_dout_14_ )
  );
  AOI22X1 _06999_ (
    .A( dbg_0.mem_data_15_ ),
    .B(_00311_),
    .C(_00514_),
    .D( dbg_0.mem_cnt_15_ ),
    .Y(_00650_)
  );
  AOI22X1 _07000_ (
    .A(1'h0),
    .B(_00582_),
    .C(_00583_),
    .D(1'h1),
    .Y(_00651_)
  );
  AOI22X1 _07001_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B(_00451_),
    .C(_00584_),
    .D(1'h0),
    .Y(_00652_)
  );
  NAND3X1 _07002_ (
    .A(_00650_),
    .B(_00651_),
    .C(_00652_),
    .Y( dbg_0.dbg_dout_15_ )
  );
  OAI21X1 _07003_ (
    .A( dbg_0.cpu_ctl_4_ ),
    .B(_00297_),
    .C( dbg_0.cpu_stat_full_0_ ),
    .Y(_00653_)
  );
  INVX1 _07004_ (
    .A(_00653_),
    .Y(_06214_)
  );
  AND2X1 _07005_ (
    .A(_00298_),
    .B(_00435_),
    .Y( dbg_0.dbg_halt_cmd )
  );
  NOR2X1 _07006_ (
    .A(_00259_),
    .B(_00439_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_wr )
  );
  OAI21X1 _07007_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_i2c_0.dbg_rd ),
    .C( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00654_)
  );
  OAI21X1 _07008_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00439_),
    .C(_00654_),
    .Y(_00166_)
  );
  AND2X1 _07009_ (
    .A(_00259_),
    .B( dbg_0.dbg_mem_en ),
    .Y( dbg_0.dbg_mem_rd )
  );
  INVX1 _07010_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00168_)
  );
  INVX1 _07011_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00169_)
  );
  INVX1 _07012_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00170_)
  );
  INVX1 _07013_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00171_)
  );
  INVX1 _07014_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00172_)
  );
  INVX1 _07015_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00173_)
  );
  INVX1 _07016_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00174_)
  );
  INVX1 _07017_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00175_)
  );
  INVX1 _07018_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00176_)
  );
  INVX1 _07019_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00177_)
  );
  INVX1 _07020_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00178_)
  );
  INVX1 _07021_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00179_)
  );
  INVX1 _07022_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00180_)
  );
  INVX1 _07023_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00181_)
  );
  INVX1 _07024_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00182_)
  );
  INVX1 _07025_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00183_)
  );
  INVX1 _07026_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00184_)
  );
  INVX1 _07027_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00185_)
  );
  INVX1 _07028_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00186_)
  );
  INVX1 _07029_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00187_)
  );
  INVX1 _07030_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00188_)
  );
  INVX1 _07031_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00189_)
  );
  INVX1 _07032_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00190_)
  );
  INVX1 _07033_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00191_)
  );
  INVX1 _07034_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00192_)
  );
  INVX1 _07035_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00193_)
  );
  INVX1 _07036_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00194_)
  );
  INVX1 _07037_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00195_)
  );
  INVX1 _07038_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00196_)
  );
  INVX1 _07039_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00197_)
  );
  INVX1 _07040_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00198_)
  );
  INVX1 _07041_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00199_)
  );
  INVX1 _07042_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00200_)
  );
  INVX1 _07043_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00201_)
  );
  INVX1 _07044_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00202_)
  );
  INVX1 _07045_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00203_)
  );
  INVX1 _07046_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00204_)
  );
  INVX1 _07047_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00205_)
  );
  INVX1 _07048_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00206_)
  );
  INVX1 _07049_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00207_)
  );
  INVX1 _07050_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00208_)
  );
  INVX1 _07051_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00209_)
  );
  INVX1 _07052_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00210_)
  );
  INVX1 _07053_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00211_)
  );
  INVX1 _07054_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00212_)
  );
  INVX1 _07055_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00213_)
  );
  INVX1 _07056_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00214_)
  );
  INVX1 _07057_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00215_)
  );
  INVX1 _07058_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00216_)
  );
  INVX1 _07059_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00217_)
  );
  INVX1 _07060_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00218_)
  );
  INVX1 _07061_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00219_)
  );
  INVX1 _07062_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00220_)
  );
  INVX1 _07063_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00221_)
  );
  INVX1 _07064_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00222_)
  );
  INVX1 _07065_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00223_)
  );
  INVX1 _07066_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00224_)
  );
  INVX1 _07067_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00225_)
  );
  INVX1 _07068_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00226_)
  );
  INVX1 _07069_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00227_)
  );
  INVX1 _07070_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00228_)
  );
  INVX1 _07071_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00229_)
  );
  INVX1 _07072_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00230_)
  );
  INVX1 _07073_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00231_)
  );
  INVX1 _07074_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00232_)
  );
  INVX1 _07075_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00233_)
  );
  DFFSR _07076_ (
    .CLK(dco_clk),
    .D(_00234_),
    .Q( dbg_0.cpu_ctl_3_ ),
    .R(_00167_),
    .S(1'h1)
  );
  DFFSR _07077_ (
    .CLK(dco_clk),
    .D(_00235_),
    .Q( dbg_0.cpu_ctl_4_ ),
    .R(1'h1),
    .S(_00168_)
  );
  DFFSR _07078_ (
    .CLK(dco_clk),
    .D(_00236_),
    .Q( dbg_0.cpu_ctl_5_ ),
    .R(_00169_),
    .S(1'h1)
  );
  DFFSR _07079_ (
    .CLK(dco_clk),
    .D(_00237_),
    .Q( clock_module_0.dbg_cpu_reset ),
    .R(_00170_),
    .S(1'h1)
  );
  DFFSR _07080_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_mem_rd ),
    .Q( dbg_0.dbg_mem_rd_dly ),
    .R(_00171_),
    .S(1'h1)
  );
  DFFSR _07081_ (
    .CLK(dco_clk),
    .D( dbg_0.mem_state_nxt_0_ ),
    .Q( dbg_0.mem_state_0_ ),
    .R(_00172_),
    .S(1'h1)
  );
  DFFSR _07082_ (
    .CLK(dco_clk),
    .D( dbg_0.mem_state_nxt_1_ ),
    .Q( dbg_0.mem_state_1_ ),
    .R(_00173_),
    .S(1'h1)
  );
  DFFSR _07083_ (
    .CLK(dco_clk),
    .D(_00166_),
    .Q( dbg_0.mem_startb ),
    .R(_00174_),
    .S(1'h1)
  );
  DFFSR _07084_ (
    .CLK(dco_clk),
    .D(_00238_),
    .Q( dbg_0.dbg_i2c_0.mem_burst ),
    .R(_00175_),
    .S(1'h1)
  );
  DFFSR _07085_ (
    .CLK(dco_clk),
    .D( dbg_0.istep ),
    .Q( dbg_0.inc_step_0_ ),
    .R(_00176_),
    .S(1'h1)
  );
  DFFSR _07086_ (
    .CLK(dco_clk),
    .D(_00132_),
    .Q( dbg_0.inc_step_1_ ),
    .R(_00177_),
    .S(1'h1)
  );
  DFFSR _07087_ (
    .CLK(dco_clk),
    .D(_00131_),
    .Q( dbg_0.dbg_rd_rdy ),
    .R(_00178_),
    .S(1'h1)
  );
  DFFSR _07088_ (
    .CLK(dco_clk),
    .D(_00149_),
    .Q( dbg_0.mem_cnt_0_ ),
    .R(_00179_),
    .S(1'h1)
  );
  DFFSR _07089_ (
    .CLK(dco_clk),
    .D(_00156_),
    .Q( dbg_0.mem_cnt_1_ ),
    .R(_00180_),
    .S(1'h1)
  );
  DFFSR _07090_ (
    .CLK(dco_clk),
    .D(_00157_),
    .Q( dbg_0.mem_cnt_2_ ),
    .R(_00181_),
    .S(1'h1)
  );
  DFFSR _07091_ (
    .CLK(dco_clk),
    .D(_00158_),
    .Q( dbg_0.mem_cnt_3_ ),
    .R(_00182_),
    .S(1'h1)
  );
  DFFSR _07092_ (
    .CLK(dco_clk),
    .D(_00159_),
    .Q( dbg_0.mem_cnt_4_ ),
    .R(_00183_),
    .S(1'h1)
  );
  DFFSR _07093_ (
    .CLK(dco_clk),
    .D(_00160_),
    .Q( dbg_0.mem_cnt_5_ ),
    .R(_00184_),
    .S(1'h1)
  );
  DFFSR _07094_ (
    .CLK(dco_clk),
    .D(_00161_),
    .Q( dbg_0.mem_cnt_6_ ),
    .R(_00185_),
    .S(1'h1)
  );
  DFFSR _07095_ (
    .CLK(dco_clk),
    .D(_00162_),
    .Q( dbg_0.mem_cnt_7_ ),
    .R(_00186_),
    .S(1'h1)
  );
  DFFSR _07096_ (
    .CLK(dco_clk),
    .D(_00163_),
    .Q( dbg_0.mem_cnt_8_ ),
    .R(_00187_),
    .S(1'h1)
  );
  DFFSR _07097_ (
    .CLK(dco_clk),
    .D(_00164_),
    .Q( dbg_0.mem_cnt_9_ ),
    .R(_00188_),
    .S(1'h1)
  );
  DFFSR _07098_ (
    .CLK(dco_clk),
    .D(_00150_),
    .Q( dbg_0.mem_cnt_10_ ),
    .R(_00189_),
    .S(1'h1)
  );
  DFFSR _07099_ (
    .CLK(dco_clk),
    .D(_00151_),
    .Q( dbg_0.mem_cnt_11_ ),
    .R(_00190_),
    .S(1'h1)
  );
  DFFSR _07100_ (
    .CLK(dco_clk),
    .D(_00152_),
    .Q( dbg_0.mem_cnt_12_ ),
    .R(_00191_),
    .S(1'h1)
  );
  DFFSR _07101_ (
    .CLK(dco_clk),
    .D(_00153_),
    .Q( dbg_0.mem_cnt_13_ ),
    .R(_00192_),
    .S(1'h1)
  );
  DFFSR _07102_ (
    .CLK(dco_clk),
    .D(_00154_),
    .Q( dbg_0.mem_cnt_14_ ),
    .R(_00193_),
    .S(1'h1)
  );
  DFFSR _07103_ (
    .CLK(dco_clk),
    .D(_00155_),
    .Q( dbg_0.mem_cnt_15_ ),
    .R(_00194_),
    .S(1'h1)
  );
  DFFSR _07104_ (
    .CLK(dco_clk),
    .D(_00133_),
    .Q( dbg_0.dbg_mem_addr_0_ ),
    .R(_00195_),
    .S(1'h1)
  );
  DFFSR _07105_ (
    .CLK(dco_clk),
    .D(_00140_),
    .Q( dbg_0.dbg_mem_addr_1_ ),
    .R(_00196_),
    .S(1'h1)
  );
  DFFSR _07106_ (
    .CLK(dco_clk),
    .D(_00141_),
    .Q( dbg_0.dbg_mem_addr_2_ ),
    .R(_00197_),
    .S(1'h1)
  );
  DFFSR _07107_ (
    .CLK(dco_clk),
    .D(_00142_),
    .Q( dbg_0.dbg_mem_addr_3_ ),
    .R(_00198_),
    .S(1'h1)
  );
  DFFSR _07108_ (
    .CLK(dco_clk),
    .D(_00143_),
    .Q( dbg_0.dbg_mem_addr_4_ ),
    .R(_00199_),
    .S(1'h1)
  );
  DFFSR _07109_ (
    .CLK(dco_clk),
    .D(_00144_),
    .Q( dbg_0.dbg_mem_addr_5_ ),
    .R(_00200_),
    .S(1'h1)
  );
  DFFSR _07110_ (
    .CLK(dco_clk),
    .D(_00145_),
    .Q( dbg_0.dbg_mem_addr_6_ ),
    .R(_00201_),
    .S(1'h1)
  );
  DFFSR _07111_ (
    .CLK(dco_clk),
    .D(_00146_),
    .Q( dbg_0.dbg_mem_addr_7_ ),
    .R(_00202_),
    .S(1'h1)
  );
  DFFSR _07112_ (
    .CLK(dco_clk),
    .D(_00147_),
    .Q( dbg_0.dbg_mem_addr_8_ ),
    .R(_00203_),
    .S(1'h1)
  );
  DFFSR _07113_ (
    .CLK(dco_clk),
    .D(_00148_),
    .Q( dbg_0.dbg_mem_addr_9_ ),
    .R(_00204_),
    .S(1'h1)
  );
  DFFSR _07114_ (
    .CLK(dco_clk),
    .D(_00134_),
    .Q( dbg_0.dbg_mem_addr_10_ ),
    .R(_00205_),
    .S(1'h1)
  );
  DFFSR _07115_ (
    .CLK(dco_clk),
    .D(_00135_),
    .Q( dbg_0.dbg_mem_addr_11_ ),
    .R(_00206_),
    .S(1'h1)
  );
  DFFSR _07116_ (
    .CLK(dco_clk),
    .D(_00136_),
    .Q( dbg_0.dbg_mem_addr_12_ ),
    .R(_00207_),
    .S(1'h1)
  );
  DFFSR _07117_ (
    .CLK(dco_clk),
    .D(_00137_),
    .Q( dbg_0.dbg_mem_addr_13_ ),
    .R(_00208_),
    .S(1'h1)
  );
  DFFSR _07118_ (
    .CLK(dco_clk),
    .D(_00138_),
    .Q( dbg_0.dbg_mem_addr_14_ ),
    .R(_00209_),
    .S(1'h1)
  );
  DFFSR _07119_ (
    .CLK(dco_clk),
    .D(_00139_),
    .Q( dbg_0.dbg_mem_addr_15_ ),
    .R(_00210_),
    .S(1'h1)
  );
  DFFSR _07120_ (
    .CLK(dco_clk),
    .D(_00239_),
    .Q( dbg_0.halt_flag ),
    .R(_00211_),
    .S(1'h1)
  );
  DFFSR _07121_ (
    .CLK(dco_clk),
    .D(_00165_),
    .Q( dbg_0.mem_start ),
    .R(_00212_),
    .S(1'h1)
  );
  DFFSR _07122_ (
    .CLK(dco_clk),
    .D(_00240_),
    .Q( dbg_0.mem_data_0_ ),
    .R(_00213_),
    .S(1'h1)
  );
  DFFSR _07123_ (
    .CLK(dco_clk),
    .D(_00241_),
    .Q( dbg_0.mem_data_1_ ),
    .R(_00214_),
    .S(1'h1)
  );
  DFFSR _07124_ (
    .CLK(dco_clk),
    .D(_00242_),
    .Q( dbg_0.mem_data_2_ ),
    .R(_00215_),
    .S(1'h1)
  );
  DFFSR _07125_ (
    .CLK(dco_clk),
    .D(_00243_),
    .Q( dbg_0.mem_data_3_ ),
    .R(_00216_),
    .S(1'h1)
  );
  DFFSR _07126_ (
    .CLK(dco_clk),
    .D(_00244_),
    .Q( dbg_0.mem_data_4_ ),
    .R(_00217_),
    .S(1'h1)
  );
  DFFSR _07127_ (
    .CLK(dco_clk),
    .D(_00245_),
    .Q( dbg_0.mem_data_5_ ),
    .R(_00218_),
    .S(1'h1)
  );
  DFFSR _07128_ (
    .CLK(dco_clk),
    .D(_00246_),
    .Q( dbg_0.mem_data_6_ ),
    .R(_00219_),
    .S(1'h1)
  );
  DFFSR _07129_ (
    .CLK(dco_clk),
    .D(_00247_),
    .Q( dbg_0.mem_data_7_ ),
    .R(_00220_),
    .S(1'h1)
  );
  DFFSR _07130_ (
    .CLK(dco_clk),
    .D(_00248_),
    .Q( dbg_0.mem_data_8_ ),
    .R(_00221_),
    .S(1'h1)
  );
  DFFSR _07131_ (
    .CLK(dco_clk),
    .D(_00249_),
    .Q( dbg_0.mem_data_9_ ),
    .R(_00222_),
    .S(1'h1)
  );
  DFFSR _07132_ (
    .CLK(dco_clk),
    .D(_00250_),
    .Q( dbg_0.mem_data_10_ ),
    .R(_00223_),
    .S(1'h1)
  );
  DFFSR _07133_ (
    .CLK(dco_clk),
    .D(_00251_),
    .Q( dbg_0.mem_data_11_ ),
    .R(_00224_),
    .S(1'h1)
  );
  DFFSR _07134_ (
    .CLK(dco_clk),
    .D(_00252_),
    .Q( dbg_0.mem_data_12_ ),
    .R(_00225_),
    .S(1'h1)
  );
  DFFSR _07135_ (
    .CLK(dco_clk),
    .D(_00253_),
    .Q( dbg_0.mem_data_13_ ),
    .R(_00226_),
    .S(1'h1)
  );
  DFFSR _07136_ (
    .CLK(dco_clk),
    .D(_00254_),
    .Q( dbg_0.mem_data_14_ ),
    .R(_00227_),
    .S(1'h1)
  );
  DFFSR _07137_ (
    .CLK(dco_clk),
    .D(_00255_),
    .Q( dbg_0.mem_data_15_ ),
    .R(_00228_),
    .S(1'h1)
  );
  DFFSR _07138_ (
    .CLK(dco_clk),
    .D(_00129_),
    .Q( dbg_0.cpu_stat_2_ ),
    .R(_00229_),
    .S(1'h1)
  );
  DFFSR _07139_ (
    .CLK(dco_clk),
    .D(_00130_),
    .Q( dbg_0.cpu_stat_3_ ),
    .R(_00230_),
    .S(1'h1)
  );
  DFFSR _07140_ (
    .CLK(dco_clk),
    .D(_00256_),
    .Q( dbg_0.mem_ctl_1_ ),
    .R(_00231_),
    .S(1'h1)
  );
  DFFSR _07141_ (
    .CLK(dco_clk),
    .D(_00257_),
    .Q( dbg_0.mem_ctl_2_ ),
    .R(_00232_),
    .S(1'h1)
  );
  DFFSR _07142_ (
    .CLK(dco_clk),
    .D(_00258_),
    .Q( dbg_0.dbg_i2c_0.mem_bw ),
    .R(_00233_),
    .S(1'h1)
  );
  INVX1 _07143_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .Y(_00741_)
  );
  INVX1 _07144_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00742_)
  );
  INVX1 _07145_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .Y(_00743_)
  );
  INVX1 _07146_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00744_)
  );
  INVX1 _07147_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .Y(_00745_)
  );
  INVX1 _07148_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00746_)
  );
  INVX1 _07149_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .Y(_00747_)
  );
  INVX1 _07150_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00748_)
  );
  INVX1 _07151_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .Y(_00749_)
  );
  INVX1 _07152_ (
    .A( dbg_0.dbg_i2c_0.dbg_bw ),
    .Y(_00750_)
  );
  INVX1 _07153_ (
    .A( dbg_0.dbg_din_15_ ),
    .Y(_00751_)
  );
  INVX1 _07154_ (
    .A( dbg_0.dbg_din_14_ ),
    .Y(_00752_)
  );
  INVX1 _07155_ (
    .A( dbg_0.dbg_din_13_ ),
    .Y(_00753_)
  );
  INVX1 _07156_ (
    .A( dbg_0.dbg_din_12_ ),
    .Y(_00754_)
  );
  INVX1 _07157_ (
    .A( dbg_0.dbg_din_11_ ),
    .Y(_00755_)
  );
  INVX1 _07158_ (
    .A( dbg_0.dbg_din_10_ ),
    .Y(_00756_)
  );
  INVX1 _07159_ (
    .A( dbg_0.dbg_din_9_ ),
    .Y(_00757_)
  );
  INVX1 _07160_ (
    .A( dbg_0.dbg_din_8_ ),
    .Y(_00758_)
  );
  INVX1 _07161_ (
    .A( dbg_0.dbg_i2c_0.scl_sync_n ),
    .Y( dbg_0.dbg_i2c_0.scl_sync )
  );
  INVX1 _07162_ (
    .A( dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .Y( dbg_0.dbg_i2c_0.sda_in_sync )
  );
  INVX1 _07163_ (
    .A( dbg_0.dbg_i2c_0.sda_in_dly ),
    .Y(_00759_)
  );
  INVX1 _07164_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00760_)
  );
  INVX1 _07165_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00761_)
  );
  INVX1 _07166_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00762_)
  );
  INVX1 _07167_ (
    .A(dbg_i2c_addr_2_),
    .Y(_00763_)
  );
  INVX1 _07168_ (
    .A(dbg_i2c_addr_3_),
    .Y(_00764_)
  );
  INVX1 _07169_ (
    .A(dbg_i2c_addr_6_),
    .Y(_00765_)
  );
  INVX1 _07170_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00766_)
  );
  INVX1 _07171_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00767_)
  );
  INVX1 _07172_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00768_)
  );
  INVX1 _07173_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00769_)
  );
  INVX1 _07174_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_wr ),
    .Y(_00770_)
  );
  INVX1 _07175_ (
    .A(dbg_i2c_scl),
    .Y( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in )
  );
  INVX1 _07176_ (
    .A(dbg_i2c_sda_in),
    .Y( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in )
  );
  INVX1 _07177_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00657_)
  );
  OR2X1 _07178_ (
    .A( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .Y(_00771_)
  );
  AND2X1 _07179_ (
    .A( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .Y(_00772_)
  );
  OAI21X1 _07180_ (
    .A( dbg_0.dbg_i2c_0.scl_sync ),
    .B(_00772_),
    .C(_00771_),
    .Y(_00773_)
  );
  INVX1 _07181_ (
    .A(_00773_),
    .Y( dbg_0.dbg_i2c_0.scl )
  );
  OR2X1 _07182_ (
    .A( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .Y(_00774_)
  );
  AND2X1 _07183_ (
    .A( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .Y(_00775_)
  );
  OAI21X1 _07184_ (
    .A( dbg_0.dbg_i2c_0.sda_in_sync ),
    .B(_00775_),
    .C(_00774_),
    .Y(_00776_)
  );
  INVX1 _07185_ (
    .A(_00776_),
    .Y( dbg_0.dbg_i2c_0.sda_in )
  );
  NAND3X1 _07186_ (
    .A( dbg_0.dbg_i2c_0.sda_in_dly ),
    .B( dbg_0.dbg_i2c_0.scl ),
    .C(_00776_),
    .Y(_00777_)
  );
  AND2X1 _07187_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00773_),
    .Y(_00778_)
  );
  NAND2X1 _07188_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00773_),
    .Y(_00779_)
  );
  NOR2X1 _07189_ (
    .A(_00741_),
    .B( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00780_)
  );
  NAND3X1 _07190_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00773_),
    .C(_00780_),
    .Y(_00781_)
  );
  AOI21X1 _07191_ (
    .A(_00761_),
    .B( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .C( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00782_)
  );
  NAND2X1 _07192_ (
    .A(_00761_),
    .B(_00782_),
    .Y(_00783_)
  );
  NOR2X1 _07193_ (
    .A(_00781_),
    .B(_00783_),
    .Y(_00784_)
  );
  INVX1 _07194_ (
    .A(_00784_),
    .Y(_00785_)
  );
  XOR2X1 _07195_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_i2c_addr_5_),
    .Y(_00786_)
  );
  NOR2X1 _07196_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_i2c_addr_1_),
    .Y(_00787_)
  );
  AND2X1 _07197_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_i2c_addr_1_),
    .Y(_00788_)
  );
  AOI21X1 _07198_ (
    .A(_00742_),
    .B(dbg_i2c_addr_6_),
    .C(_00786_),
    .Y(_00789_)
  );
  AOI22X1 _07199_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00764_),
    .C(dbg_i2c_addr_4_),
    .D(_00744_),
    .Y(_00790_)
  );
  AOI22X1 _07200_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00763_),
    .C(_00765_),
    .D( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00791_)
  );
  NAND3X1 _07201_ (
    .A(_00789_),
    .B(_00790_),
    .C(_00791_),
    .Y(_00792_)
  );
  XNOR2X1 _07202_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(dbg_i2c_addr_0_),
    .Y(_00793_)
  );
  OAI21X1 _07203_ (
    .A(_00787_),
    .B(_00788_),
    .C(_00793_),
    .Y(_00794_)
  );
  AOI22X1 _07204_ (
    .A(_00746_),
    .B(dbg_i2c_addr_2_),
    .C(dbg_i2c_addr_3_),
    .D(_00745_),
    .Y(_00795_)
  );
  OAI21X1 _07205_ (
    .A(_00744_),
    .B(dbg_i2c_addr_4_),
    .C(_00795_),
    .Y(_00796_)
  );
  NOR3X1 _07206_ (
    .A(_00792_),
    .B(_00794_),
    .C(_00796_),
    .Y(_00797_)
  );
  NOR2X1 _07207_ (
    .A(_00785_),
    .B(_00797_),
    .Y(_00798_)
  );
  NAND3X1 _07208_ (
    .A(_00759_),
    .B( dbg_0.dbg_i2c_0.scl ),
    .C( dbg_0.dbg_i2c_0.sda_in ),
    .Y(_00799_)
  );
  NAND2X1 _07209_ (
    .A( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .B(_00799_),
    .Y(_00800_)
  );
  OAI21X1 _07210_ (
    .A(_00798_),
    .B(_00800_),
    .C(_00777_),
    .Y(_00740_)
  );
  NAND3X1 _07211_ (
    .A( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .B(_00777_),
    .C(_00799_),
    .Y(_00801_)
  );
  NAND2X1 _07212_ (
    .A(_00760_),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00802_)
  );
  OR2X1 _07213_ (
    .A(_00762_),
    .B(_00802_),
    .Y(_00803_)
  );
  NOR3X1 _07214_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .C(_00762_),
    .Y(_00804_)
  );
  NAND3X1 _07215_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00773_),
    .C(_00804_),
    .Y(_00805_)
  );
  OR2X1 _07216_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00805_),
    .Y(_00806_)
  );
  OAI22X1 _07217_ (
    .A(_00779_),
    .B(_00803_),
    .C(_00805_),
    .D( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .Y(_00807_)
  );
  NOR2X1 _07218_ (
    .A(_00801_),
    .B(_00807_),
    .Y(_00808_)
  );
  NOR2X1 _07219_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00809_)
  );
  NOR2X1 _07220_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00773_),
    .Y( dbg_0.dbg_i2c_0.scl_re )
  );
  NAND3X1 _07221_ (
    .A(_00761_),
    .B( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .C( dbg_0.dbg_i2c_0.scl_re ),
    .Y(_00810_)
  );
  OR2X1 _07222_ (
    .A(_00809_),
    .B(_00810_),
    .Y(_00811_)
  );
  AND2X1 _07223_ (
    .A(_00808_),
    .B(_00811_),
    .Y(_00812_)
  );
  OR2X1 _07224_ (
    .A(_00749_),
    .B(_00805_),
    .Y(_00813_)
  );
  NOR2X1 _07225_ (
    .A(_00760_),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00814_)
  );
  NAND2X1 _07226_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .B( dbg_0.dbg_i2c_0.sda_in ),
    .Y(_00815_)
  );
  OAI21X1 _07227_ (
    .A(_00779_),
    .B(_00815_),
    .C(_00814_),
    .Y(_00816_)
  );
  OAI21X1 _07228_ (
    .A(_00749_),
    .B(_00805_),
    .C(_00816_),
    .Y(_00817_)
  );
  AOI21X1 _07229_ (
    .A(_00813_),
    .B(_00816_),
    .C(_00801_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ )
  );
  NOR2X1 _07230_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00818_)
  );
  NAND2X1 _07231_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00742_),
    .Y(_00819_)
  );
  NOR2X1 _07232_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00820_)
  );
  NAND3X1 _07233_ (
    .A(_00743_),
    .B(_00744_),
    .C(_00820_),
    .Y(_00821_)
  );
  NOR2X1 _07234_ (
    .A(_00819_),
    .B(_00821_),
    .Y(_00822_)
  );
  NAND3X1 _07235_ (
    .A(_00749_),
    .B(_00818_),
    .C(_00822_),
    .Y(_00823_)
  );
  NAND3X1 _07236_ (
    .A(_00778_),
    .B( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ),
    .C(_00823_),
    .Y(_00824_)
  );
  NAND2X1 _07237_ (
    .A( dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .B(_00782_),
    .Y(_00825_)
  );
  NAND3X1 _07238_ (
    .A(_00812_),
    .B(_00824_),
    .C(_00825_),
    .Y(_00826_)
  );
  NAND3X1 _07239_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00766_),
    .C(_00767_),
    .Y(_00827_)
  );
  MUX2X1 _07240_ (
    .A( dbg_0.dbg_dout_7_ ),
    .B( dbg_0.dbg_dout_15_ ),
    .S(_00827_),
    .Y(_00828_)
  );
  MUX2X1 _07241_ (
    .A(_00742_),
    .B(_00828_),
    .S(_00811_),
    .Y(_00829_)
  );
  NAND2X1 _07242_ (
    .A(_00808_),
    .B(_00829_),
    .Y(_00830_)
  );
  MUX2X1 _07243_ (
    .A(_00830_),
    .B(_00741_),
    .S(_00826_),
    .Y(_00739_)
  );
  MUX2X1 _07244_ (
    .A( dbg_0.dbg_dout_6_ ),
    .B( dbg_0.dbg_dout_14_ ),
    .S(_00827_),
    .Y(_00831_)
  );
  MUX2X1 _07245_ (
    .A(_00743_),
    .B(_00831_),
    .S(_00811_),
    .Y(_00832_)
  );
  NAND2X1 _07246_ (
    .A(_00808_),
    .B(_00832_),
    .Y(_00833_)
  );
  MUX2X1 _07247_ (
    .A(_00833_),
    .B(_00742_),
    .S(_00826_),
    .Y(_00738_)
  );
  MUX2X1 _07248_ (
    .A( dbg_0.dbg_dout_5_ ),
    .B( dbg_0.dbg_dout_13_ ),
    .S(_00827_),
    .Y(_00834_)
  );
  MUX2X1 _07249_ (
    .A(_00744_),
    .B(_00834_),
    .S(_00811_),
    .Y(_00835_)
  );
  NAND2X1 _07250_ (
    .A(_00808_),
    .B(_00835_),
    .Y(_00836_)
  );
  MUX2X1 _07251_ (
    .A(_00836_),
    .B(_00743_),
    .S(_00826_),
    .Y(_00737_)
  );
  MUX2X1 _07252_ (
    .A( dbg_0.dbg_dout_4_ ),
    .B( dbg_0.dbg_dout_12_ ),
    .S(_00827_),
    .Y(_00837_)
  );
  MUX2X1 _07253_ (
    .A(_00745_),
    .B(_00837_),
    .S(_00811_),
    .Y(_00838_)
  );
  NAND2X1 _07254_ (
    .A(_00808_),
    .B(_00838_),
    .Y(_00839_)
  );
  MUX2X1 _07255_ (
    .A(_00839_),
    .B(_00744_),
    .S(_00826_),
    .Y(_00736_)
  );
  MUX2X1 _07256_ (
    .A( dbg_0.dbg_dout_3_ ),
    .B( dbg_0.dbg_dout_11_ ),
    .S(_00827_),
    .Y(_00840_)
  );
  MUX2X1 _07257_ (
    .A(_00746_),
    .B(_00840_),
    .S(_00811_),
    .Y(_00841_)
  );
  NAND2X1 _07258_ (
    .A(_00808_),
    .B(_00841_),
    .Y(_00842_)
  );
  MUX2X1 _07259_ (
    .A(_00842_),
    .B(_00745_),
    .S(_00826_),
    .Y(_00735_)
  );
  MUX2X1 _07260_ (
    .A( dbg_0.dbg_dout_2_ ),
    .B( dbg_0.dbg_dout_10_ ),
    .S(_00827_),
    .Y(_00843_)
  );
  MUX2X1 _07261_ (
    .A(_00747_),
    .B(_00843_),
    .S(_00811_),
    .Y(_00844_)
  );
  NAND2X1 _07262_ (
    .A(_00808_),
    .B(_00844_),
    .Y(_00845_)
  );
  MUX2X1 _07263_ (
    .A(_00845_),
    .B(_00746_),
    .S(_00826_),
    .Y(_00734_)
  );
  MUX2X1 _07264_ (
    .A( dbg_0.dbg_dout_1_ ),
    .B( dbg_0.dbg_dout_9_ ),
    .S(_00827_),
    .Y(_00846_)
  );
  MUX2X1 _07265_ (
    .A(_00748_),
    .B(_00846_),
    .S(_00811_),
    .Y(_00847_)
  );
  NAND2X1 _07266_ (
    .A(_00808_),
    .B(_00847_),
    .Y(_00848_)
  );
  MUX2X1 _07267_ (
    .A(_00848_),
    .B(_00747_),
    .S(_00826_),
    .Y(_00733_)
  );
  NAND2X1 _07268_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00810_),
    .Y(_00849_)
  );
  MUX2X1 _07269_ (
    .A( dbg_0.dbg_dout_0_ ),
    .B( dbg_0.dbg_dout_8_ ),
    .S(_00827_),
    .Y(_00850_)
  );
  OAI21X1 _07270_ (
    .A(_00811_),
    .B(_00850_),
    .C(_00849_),
    .Y(_00851_)
  );
  NAND2X1 _07271_ (
    .A(_00808_),
    .B(_00851_),
    .Y(_00852_)
  );
  MUX2X1 _07272_ (
    .A(_00852_),
    .B(_00748_),
    .S(_00826_),
    .Y(_00732_)
  );
  OR2X1 _07273_ (
    .A(_00776_),
    .B(_00825_),
    .Y(_00853_)
  );
  AND2X1 _07274_ (
    .A(_00812_),
    .B(_00853_),
    .Y(_00854_)
  );
  OAI21X1 _07275_ (
    .A(_00749_),
    .B(_00826_),
    .C(_00854_),
    .Y(_00731_)
  );
  NAND2X1 _07276_ (
    .A(_06215_),
    .B(_00779_),
    .Y(_00855_)
  );
  AND2X1 _07277_ (
    .A(_00784_),
    .B(_00797_),
    .Y(_00856_)
  );
  NOR2X1 _07278_ (
    .A(_00781_),
    .B(_00802_),
    .Y(_00857_)
  );
  OAI21X1 _07279_ (
    .A(_00760_),
    .B(_00761_),
    .C( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00858_)
  );
  OAI22X1 _07280_ (
    .A(_00781_),
    .B(_00802_),
    .C(_00858_),
    .D(_00778_),
    .Y(_00859_)
  );
  NAND2X1 _07281_ (
    .A(_00778_),
    .B(_00814_),
    .Y(_00860_)
  );
  NOR2X1 _07282_ (
    .A(_00823_),
    .B(_00860_),
    .Y(_00861_)
  );
  OR2X1 _07283_ (
    .A(_00823_),
    .B(_00860_),
    .Y(_00862_)
  );
  NOR3X1 _07284_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .B(_00823_),
    .C(_00860_),
    .Y(_00863_)
  );
  NOR3X1 _07285_ (
    .A(_00856_),
    .B(_00859_),
    .C(_00863_),
    .Y(_00864_)
  );
  NOR2X1 _07286_ (
    .A(_00801_),
    .B(_00864_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_0_ )
  );
  NOR3X1 _07287_ (
    .A(_00801_),
    .B(_00817_),
    .C(_00864_),
    .Y(_00865_)
  );
  OAI21X1 _07288_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00824_),
    .C(_00778_),
    .Y(_00866_)
  );
  OAI21X1 _07289_ (
    .A(_00865_),
    .B(_00866_),
    .C(_00855_),
    .Y(_00730_)
  );
  NOR2X1 _07290_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00867_)
  );
  AND2X1 _07291_ (
    .A(_00767_),
    .B(_00867_),
    .Y(_00868_)
  );
  AND2X1 _07292_ (
    .A(_00857_),
    .B(_00868_),
    .Y(_00869_)
  );
  NAND2X1 _07293_ (
    .A(_00857_),
    .B(_00868_),
    .Y(_00870_)
  );
  NOR2X1 _07294_ (
    .A(_00768_),
    .B(_00769_),
    .Y(_00871_)
  );
  NAND2X1 _07295_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00872_)
  );
  AOI21X1 _07296_ (
    .A( dbg_0.dbg_i2c_0.dbg_bw ),
    .B(_00768_),
    .C(_00871_),
    .Y(_00873_)
  );
  NAND2X1 _07297_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00869_),
    .Y(_00874_)
  );
  OAI21X1 _07298_ (
    .A(_00869_),
    .B(_00873_),
    .C(_00874_),
    .Y(_00729_)
  );
  NOR2X1 _07299_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00869_),
    .Y(_00875_)
  );
  NAND2X1 _07300_ (
    .A(_00768_),
    .B(_00870_),
    .Y(_00876_)
  );
  AOI22X1 _07301_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00869_),
    .C(_00875_),
    .D( dbg_0.dbg_addr_5_ ),
    .Y(_00877_)
  );
  INVX1 _07302_ (
    .A(_00877_),
    .Y(_00728_)
  );
  AOI22X1 _07303_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00869_),
    .C(_00875_),
    .D( dbg_0.dbg_addr_4_ ),
    .Y(_00878_)
  );
  INVX1 _07304_ (
    .A(_00878_),
    .Y(_00727_)
  );
  AOI22X1 _07305_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00869_),
    .C(_00875_),
    .D( dbg_0.dbg_addr_3_ ),
    .Y(_00879_)
  );
  INVX1 _07306_ (
    .A(_00879_),
    .Y(_00726_)
  );
  OAI22X1 _07307_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(_00870_),
    .C(_00876_),
    .D( dbg_0.dbg_addr_2_ ),
    .Y(_00880_)
  );
  INVX1 _07308_ (
    .A(_00880_),
    .Y(_00725_)
  );
  OAI22X1 _07309_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(_00870_),
    .C(_00876_),
    .D( dbg_0.dbg_addr_1_ ),
    .Y(_00881_)
  );
  INVX1 _07310_ (
    .A(_00881_),
    .Y(_00724_)
  );
  AOI22X1 _07311_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00869_),
    .C(_00875_),
    .D( dbg_0.dbg_addr_0_ ),
    .Y(_00882_)
  );
  INVX1 _07312_ (
    .A(_00882_),
    .Y(_00723_)
  );
  NAND2X1 _07313_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00867_),
    .Y(_00883_)
  );
  NAND3X1 _07314_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00857_),
    .C(_00867_),
    .Y(_00884_)
  );
  MUX2X1 _07315_ (
    .A( dbg_0.dbg_din_7_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .S(_00884_),
    .Y(_00885_)
  );
  INVX1 _07316_ (
    .A(_00885_),
    .Y(_00722_)
  );
  MUX2X1 _07317_ (
    .A( dbg_0.dbg_din_6_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .S(_00884_),
    .Y(_00886_)
  );
  INVX1 _07318_ (
    .A(_00886_),
    .Y(_00721_)
  );
  MUX2X1 _07319_ (
    .A( dbg_0.dbg_din_5_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .S(_00884_),
    .Y(_00887_)
  );
  INVX1 _07320_ (
    .A(_00887_),
    .Y(_00720_)
  );
  MUX2X1 _07321_ (
    .A( dbg_0.dbg_din_4_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .S(_00884_),
    .Y(_00888_)
  );
  INVX1 _07322_ (
    .A(_00888_),
    .Y(_00719_)
  );
  MUX2X1 _07323_ (
    .A( dbg_0.dbg_din_3_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .S(_00884_),
    .Y(_00889_)
  );
  INVX1 _07324_ (
    .A(_00889_),
    .Y(_00718_)
  );
  MUX2X1 _07325_ (
    .A( dbg_0.dbg_din_2_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .S(_00884_),
    .Y(_00890_)
  );
  INVX1 _07326_ (
    .A(_00890_),
    .Y(_00717_)
  );
  MUX2X1 _07327_ (
    .A( dbg_0.dbg_din_1_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .S(_00884_),
    .Y(_00891_)
  );
  INVX1 _07328_ (
    .A(_00891_),
    .Y(_00716_)
  );
  MUX2X1 _07329_ (
    .A( dbg_0.dbg_din_0_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .S(_00884_),
    .Y(_00892_)
  );
  INVX1 _07330_ (
    .A(_00892_),
    .Y(_00715_)
  );
  OR2X1 _07331_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00766_),
    .Y(_00893_)
  );
  NOR2X1 _07332_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00893_),
    .Y(_00894_)
  );
  INVX1 _07333_ (
    .A(_00894_),
    .Y(_00895_)
  );
  NAND2X1 _07334_ (
    .A(_00857_),
    .B(_00894_),
    .Y(_00896_)
  );
  OAI21X1 _07335_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00896_),
    .C(_00884_),
    .Y(_00897_)
  );
  AOI21X1 _07336_ (
    .A(_00751_),
    .B(_00896_),
    .C(_00897_),
    .Y(_00714_)
  );
  OAI21X1 _07337_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00896_),
    .C(_00884_),
    .Y(_00898_)
  );
  AOI21X1 _07338_ (
    .A(_00752_),
    .B(_00896_),
    .C(_00898_),
    .Y(_00713_)
  );
  OAI21X1 _07339_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00896_),
    .C(_00884_),
    .Y(_00899_)
  );
  AOI21X1 _07340_ (
    .A(_00753_),
    .B(_00896_),
    .C(_00899_),
    .Y(_00712_)
  );
  NAND2X1 _07341_ (
    .A(_00884_),
    .B(_00896_),
    .Y(_00900_)
  );
  OAI22X1 _07342_ (
    .A(_00745_),
    .B(_00896_),
    .C(_00900_),
    .D(_00754_),
    .Y(_00711_)
  );
  OAI22X1 _07343_ (
    .A(_00746_),
    .B(_00896_),
    .C(_00900_),
    .D(_00755_),
    .Y(_00710_)
  );
  OAI22X1 _07344_ (
    .A(_00747_),
    .B(_00896_),
    .C(_00900_),
    .D(_00756_),
    .Y(_00709_)
  );
  OAI22X1 _07345_ (
    .A(_00748_),
    .B(_00896_),
    .C(_00900_),
    .D(_00757_),
    .Y(_00708_)
  );
  OAI22X1 _07346_ (
    .A(_00749_),
    .B(_00896_),
    .C(_00900_),
    .D(_00758_),
    .Y(_00707_)
  );
  AOI21X1 _07347_ (
    .A(_00802_),
    .B(_00806_),
    .C(_00801_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_1_ )
  );
  MUX2X1 _07348_ (
    .A(_00896_),
    .B(_00884_),
    .S(_00873_),
    .Y(_00656_)
  );
  NAND2X1 _07349_ (
    .A(_00742_),
    .B(_00869_),
    .Y(_00901_)
  );
  OR2X1 _07350_ (
    .A(_00768_),
    .B(_00827_),
    .Y(_00902_)
  );
  NOR2X1 _07351_ (
    .A(_00862_),
    .B(_00902_),
    .Y(_00903_)
  );
  OR2X1 _07352_ (
    .A(_00767_),
    .B(_00893_),
    .Y(_00904_)
  );
  NOR2X1 _07353_ (
    .A(_00862_),
    .B(_00904_),
    .Y(_00905_)
  );
  AOI22X1 _07354_ (
    .A(_00769_),
    .B(_00903_),
    .C(_00905_),
    .D(_00871_),
    .Y(_00906_)
  );
  OAI21X1 _07355_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00901_),
    .C(_00906_),
    .Y(_00655_)
  );
  AOI21X1 _07356_ (
    .A(_00861_),
    .B(_00872_),
    .C(_00904_),
    .Y(_00907_)
  );
  NOR2X1 _07357_ (
    .A(_00903_),
    .B(_00907_),
    .Y(_00908_)
  );
  OR2X1 _07358_ (
    .A(_00768_),
    .B( dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00909_)
  );
  OAI21X1 _07359_ (
    .A(_00769_),
    .B(_00909_),
    .C(_00857_),
    .Y(_00910_)
  );
  AOI21X1 _07360_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_i2c_0.mem_burst_end ),
    .C(_00883_),
    .Y(_00911_)
  );
  OAI21X1 _07361_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B( dbg_0.dbg_i2c_0.mem_burst_wr ),
    .C(_00868_),
    .Y(_00912_)
  );
  AOI21X1 _07362_ (
    .A(_00910_),
    .B(_00911_),
    .C(_00869_),
    .Y(_00913_)
  );
  OAI21X1 _07363_ (
    .A(_00896_),
    .B(_00909_),
    .C(_00912_),
    .Y(_00914_)
  );
  INVX1 _07364_ (
    .A(_00914_),
    .Y(_00915_)
  );
  NAND3X1 _07365_ (
    .A(_00908_),
    .B(_00913_),
    .C(_00915_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_0_ )
  );
  NAND2X1 _07366_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(_00868_),
    .Y(_00916_)
  );
  OAI21X1 _07367_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00870_),
    .C(_00916_),
    .Y(_00917_)
  );
  OAI21X1 _07368_ (
    .A(_00750_),
    .B( dbg_0.dbg_i2c_0.mem_burst ),
    .C(_00911_),
    .Y(_00918_)
  );
  OAI22X1 _07369_ (
    .A(_00857_),
    .B(_00895_),
    .C(_00910_),
    .D(_00918_),
    .Y(_00919_)
  );
  AOI21X1 _07370_ (
    .A(_00770_),
    .B(_00917_),
    .C(_00919_),
    .Y(_00920_)
  );
  NAND2X1 _07371_ (
    .A(_00908_),
    .B(_00920_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_1_ )
  );
  NAND2X1 _07372_ (
    .A(_00873_),
    .B(_00905_),
    .Y(_00921_)
  );
  OAI21X1 _07373_ (
    .A(_00827_),
    .B(_00861_),
    .C(_00921_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_2_ )
  );
  INVX1 _07374_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00658_)
  );
  INVX1 _07375_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00659_)
  );
  INVX1 _07376_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00660_)
  );
  INVX1 _07377_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00661_)
  );
  INVX1 _07378_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00662_)
  );
  INVX1 _07379_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00663_)
  );
  INVX1 _07380_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00664_)
  );
  INVX1 _07381_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00665_)
  );
  INVX1 _07382_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00666_)
  );
  INVX1 _07383_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00667_)
  );
  INVX1 _07384_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00668_)
  );
  INVX1 _07385_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00669_)
  );
  INVX1 _07386_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00670_)
  );
  INVX1 _07387_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00671_)
  );
  INVX1 _07388_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00672_)
  );
  INVX1 _07389_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00673_)
  );
  INVX1 _07390_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00674_)
  );
  INVX1 _07391_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00675_)
  );
  INVX1 _07392_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00676_)
  );
  INVX1 _07393_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00677_)
  );
  INVX1 _07394_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00678_)
  );
  INVX1 _07395_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00679_)
  );
  INVX1 _07396_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00680_)
  );
  INVX1 _07397_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00681_)
  );
  INVX1 _07398_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00682_)
  );
  INVX1 _07399_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00683_)
  );
  INVX1 _07400_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00684_)
  );
  INVX1 _07401_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00685_)
  );
  INVX1 _07402_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00686_)
  );
  INVX1 _07403_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00687_)
  );
  INVX1 _07404_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00688_)
  );
  INVX1 _07405_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00689_)
  );
  INVX1 _07406_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00690_)
  );
  INVX1 _07407_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00691_)
  );
  INVX1 _07408_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00692_)
  );
  INVX1 _07409_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00693_)
  );
  INVX1 _07410_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00694_)
  );
  INVX1 _07411_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00695_)
  );
  INVX1 _07412_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00696_)
  );
  INVX1 _07413_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00697_)
  );
  INVX1 _07414_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00698_)
  );
  INVX1 _07415_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00699_)
  );
  INVX1 _07416_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00700_)
  );
  INVX1 _07417_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00701_)
  );
  INVX1 _07418_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00702_)
  );
  INVX1 _07419_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00703_)
  );
  INVX1 _07420_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00704_)
  );
  INVX1 _07421_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00705_)
  );
  INVX1 _07422_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00706_)
  );
  DFFSR _07423_ (
    .CLK(dco_clk),
    .D(_00655_),
    .Q( dbg_0.dbg_i2c_0.dbg_rd ),
    .R(_00657_),
    .S(1'h1)
  );
  DFFSR _07424_ (
    .CLK(dco_clk),
    .D(_00656_),
    .Q( dbg_0.dbg_i2c_0.dbg_wr ),
    .R(_00658_),
    .S(1'h1)
  );
  DFFSR _07425_ (
    .CLK(dco_clk),
    .D(_00707_),
    .Q( dbg_0.dbg_din_8_ ),
    .R(_00659_),
    .S(1'h1)
  );
  DFFSR _07426_ (
    .CLK(dco_clk),
    .D(_00708_),
    .Q( dbg_0.dbg_din_9_ ),
    .R(_00660_),
    .S(1'h1)
  );
  DFFSR _07427_ (
    .CLK(dco_clk),
    .D(_00709_),
    .Q( dbg_0.dbg_din_10_ ),
    .R(_00661_),
    .S(1'h1)
  );
  DFFSR _07428_ (
    .CLK(dco_clk),
    .D(_00710_),
    .Q( dbg_0.dbg_din_11_ ),
    .R(_00662_),
    .S(1'h1)
  );
  DFFSR _07429_ (
    .CLK(dco_clk),
    .D(_00711_),
    .Q( dbg_0.dbg_din_12_ ),
    .R(_00663_),
    .S(1'h1)
  );
  DFFSR _07430_ (
    .CLK(dco_clk),
    .D(_00712_),
    .Q( dbg_0.dbg_din_13_ ),
    .R(_00664_),
    .S(1'h1)
  );
  DFFSR _07431_ (
    .CLK(dco_clk),
    .D(_00713_),
    .Q( dbg_0.dbg_din_14_ ),
    .R(_00665_),
    .S(1'h1)
  );
  DFFSR _07432_ (
    .CLK(dco_clk),
    .D(_00714_),
    .Q( dbg_0.dbg_din_15_ ),
    .R(_00666_),
    .S(1'h1)
  );
  DFFSR _07433_ (
    .CLK(dco_clk),
    .D(_00715_),
    .Q( dbg_0.dbg_din_0_ ),
    .R(_00667_),
    .S(1'h1)
  );
  DFFSR _07434_ (
    .CLK(dco_clk),
    .D(_00716_),
    .Q( dbg_0.dbg_din_1_ ),
    .R(_00668_),
    .S(1'h1)
  );
  DFFSR _07435_ (
    .CLK(dco_clk),
    .D(_00717_),
    .Q( dbg_0.dbg_din_2_ ),
    .R(_00669_),
    .S(1'h1)
  );
  DFFSR _07436_ (
    .CLK(dco_clk),
    .D(_00718_),
    .Q( dbg_0.dbg_din_3_ ),
    .R(_00670_),
    .S(1'h1)
  );
  DFFSR _07437_ (
    .CLK(dco_clk),
    .D(_00719_),
    .Q( dbg_0.dbg_din_4_ ),
    .R(_00671_),
    .S(1'h1)
  );
  DFFSR _07438_ (
    .CLK(dco_clk),
    .D(_00720_),
    .Q( dbg_0.dbg_din_5_ ),
    .R(_00672_),
    .S(1'h1)
  );
  DFFSR _07439_ (
    .CLK(dco_clk),
    .D(_00721_),
    .Q( dbg_0.dbg_din_6_ ),
    .R(_00673_),
    .S(1'h1)
  );
  DFFSR _07440_ (
    .CLK(dco_clk),
    .D(_00722_),
    .Q( dbg_0.dbg_din_7_ ),
    .R(_00674_),
    .S(1'h1)
  );
  DFFSR _07441_ (
    .CLK(dco_clk),
    .D(_00723_),
    .Q( dbg_0.dbg_addr_0_ ),
    .R(_00675_),
    .S(1'h1)
  );
  DFFSR _07442_ (
    .CLK(dco_clk),
    .D(_00724_),
    .Q( dbg_0.dbg_addr_1_ ),
    .R(_00676_),
    .S(1'h1)
  );
  DFFSR _07443_ (
    .CLK(dco_clk),
    .D(_00725_),
    .Q( dbg_0.dbg_addr_2_ ),
    .R(_00677_),
    .S(1'h1)
  );
  DFFSR _07444_ (
    .CLK(dco_clk),
    .D(_00726_),
    .Q( dbg_0.dbg_addr_3_ ),
    .R(_00678_),
    .S(1'h1)
  );
  DFFSR _07445_ (
    .CLK(dco_clk),
    .D(_00727_),
    .Q( dbg_0.dbg_addr_4_ ),
    .R(_00679_),
    .S(1'h1)
  );
  DFFSR _07446_ (
    .CLK(dco_clk),
    .D(_00728_),
    .Q( dbg_0.dbg_addr_5_ ),
    .R(_00680_),
    .S(1'h1)
  );
  DFFSR _07447_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_0_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .R(_00681_),
    .S(1'h1)
  );
  DFFSR _07448_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_1_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .R(_00682_),
    .S(1'h1)
  );
  DFFSR _07449_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_2_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .R(_00683_),
    .S(1'h1)
  );
  DFFSR _07450_ (
    .CLK(dco_clk),
    .D(_00729_),
    .Q( dbg_0.dbg_i2c_0.dbg_bw ),
    .R(_00684_),
    .S(1'h1)
  );
  DFFSR _07451_ (
    .CLK(dco_clk),
    .D(_00730_),
    .Q(_06215_),
    .R(1'h1),
    .S(_00685_)
  );
  DFFSR _07452_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_0_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .R(_00686_),
    .S(1'h1)
  );
  DFFSR _07453_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_1_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .R(_00687_),
    .S(1'h1)
  );
  DFFSR _07454_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .R(_00688_),
    .S(1'h1)
  );
  DFFSR _07455_ (
    .CLK(dco_clk),
    .D(_00731_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .R(1'h1),
    .S(_00689_)
  );
  DFFSR _07456_ (
    .CLK(dco_clk),
    .D(_00732_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .R(_00690_),
    .S(1'h1)
  );
  DFFSR _07457_ (
    .CLK(dco_clk),
    .D(_00733_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .R(_00691_),
    .S(1'h1)
  );
  DFFSR _07458_ (
    .CLK(dco_clk),
    .D(_00734_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .R(_00692_),
    .S(1'h1)
  );
  DFFSR _07459_ (
    .CLK(dco_clk),
    .D(_00735_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .R(_00693_),
    .S(1'h1)
  );
  DFFSR _07460_ (
    .CLK(dco_clk),
    .D(_00736_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .R(_00694_),
    .S(1'h1)
  );
  DFFSR _07461_ (
    .CLK(dco_clk),
    .D(_00737_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .R(_00695_),
    .S(1'h1)
  );
  DFFSR _07462_ (
    .CLK(dco_clk),
    .D(_00738_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .R(_00696_),
    .S(1'h1)
  );
  DFFSR _07463_ (
    .CLK(dco_clk),
    .D(_00739_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .R(_00697_),
    .S(1'h1)
  );
  DFFSR _07464_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_re ),
    .Q( dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .R(_00698_),
    .S(1'h1)
  );
  DFFSR _07465_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .R(_00699_),
    .S(1'h1)
  );
  DFFSR _07466_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl ),
    .Q( dbg_0.dbg_i2c_0.scl_dly ),
    .R(1'h1),
    .S(_00700_)
  );
  DFFSR _07467_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in ),
    .Q( dbg_0.dbg_i2c_0.sda_in_dly ),
    .R(1'h1),
    .S(_00701_)
  );
  DFFSR _07468_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in_sync ),
    .Q( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .R(1'h1),
    .S(_00702_)
  );
  DFFSR _07469_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Q( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .R(1'h1),
    .S(_00703_)
  );
  DFFSR _07470_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_sync ),
    .Q( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .R(1'h1),
    .S(_00704_)
  );
  DFFSR _07471_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .R(1'h1),
    .S(_00705_)
  );
  DFFSR _07472_ (
    .CLK(dco_clk),
    .D(_00740_),
    .Q( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .R(_00706_),
    .S(1'h1)
  );
  INVX1 _07473_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00922_)
  );
  INVX1 _07474_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00923_)
  );
  DFFSR _07475_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ),
    .Q( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .R(_00922_),
    .S(1'h1)
  );
  DFFSR _07476_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_sync_n ),
    .R(_00923_),
    .S(1'h1)
  );
  INVX1 _07477_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00924_)
  );
  INVX1 _07478_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00925_)
  );
  DFFSR _07479_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ),
    .Q( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .R(_00924_),
    .S(1'h1)
  );
  DFFSR _07480_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .Q( dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .R(_00925_),
    .S(1'h1)
  );
  INVX1 _07481_ (
    .A( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_00996_)
  );
  INVX1 _07482_ (
    .A( execution_unit_0.mdb_in_buf_15_ ),
    .Y(_00997_)
  );
  INVX1 _07483_ (
    .A( execution_unit_0.mdb_in_buf_14_ ),
    .Y(_00998_)
  );
  INVX1 _07484_ (
    .A( execution_unit_0.mdb_in_buf_13_ ),
    .Y(_00999_)
  );
  INVX1 _07485_ (
    .A( execution_unit_0.mdb_in_buf_12_ ),
    .Y(_01000_)
  );
  INVX1 _07486_ (
    .A( execution_unit_0.mdb_in_buf_11_ ),
    .Y(_01001_)
  );
  INVX1 _07487_ (
    .A( execution_unit_0.mdb_in_buf_10_ ),
    .Y(_01002_)
  );
  INVX1 _07488_ (
    .A( execution_unit_0.mdb_in_buf_9_ ),
    .Y(_01003_)
  );
  INVX1 _07489_ (
    .A( execution_unit_0.mdb_in_buf_8_ ),
    .Y(_01004_)
  );
  INVX1 _07490_ (
    .A( execution_unit_0.mdb_out_nxt_15_ ),
    .Y(_01005_)
  );
  INVX1 _07491_ (
    .A( execution_unit_0.mdb_out_nxt_14_ ),
    .Y(_01006_)
  );
  INVX1 _07492_ (
    .A( execution_unit_0.mdb_out_nxt_13_ ),
    .Y(_01007_)
  );
  INVX1 _07493_ (
    .A( execution_unit_0.mdb_out_nxt_12_ ),
    .Y(_01008_)
  );
  INVX1 _07494_ (
    .A( execution_unit_0.mdb_out_nxt_11_ ),
    .Y(_01009_)
  );
  INVX1 _07495_ (
    .A( execution_unit_0.mdb_out_nxt_10_ ),
    .Y(_01010_)
  );
  INVX1 _07496_ (
    .A( execution_unit_0.mdb_out_nxt_9_ ),
    .Y(_01011_)
  );
  INVX1 _07497_ (
    .A( execution_unit_0.mdb_out_nxt_8_ ),
    .Y(_01012_)
  );
  INVX1 _07498_ (
    .A( execution_unit_0.e_state_0_ ),
    .Y(_01013_)
  );
  INVX1 _07499_ (
    .A( execution_unit_0.e_state_2_ ),
    .Y(_01014_)
  );
  INVX1 _07500_ (
    .A( execution_unit_0.e_state_3_ ),
    .Y(_01015_)
  );
  INVX1 _07501_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01016_)
  );
  INVX1 _07502_ (
    .A( execution_unit_0.inst_as_5_ ),
    .Y(_01017_)
  );
  INVX1 _07503_ (
    .A( dbg_0.dbg_reg_din_0_ ),
    .Y(_01018_)
  );
  INVX1 _07504_ (
    .A( dbg_0.dbg_reg_din_1_ ),
    .Y(_01019_)
  );
  INVX1 _07505_ (
    .A( dbg_0.dbg_reg_din_2_ ),
    .Y(_01020_)
  );
  INVX1 _07506_ (
    .A( dbg_0.dbg_reg_din_3_ ),
    .Y(_01021_)
  );
  INVX1 _07507_ (
    .A( dbg_0.dbg_reg_din_4_ ),
    .Y(_01022_)
  );
  INVX1 _07508_ (
    .A( dbg_0.dbg_reg_din_5_ ),
    .Y(_01023_)
  );
  INVX1 _07509_ (
    .A( dbg_0.dbg_reg_din_6_ ),
    .Y(_01024_)
  );
  INVX1 _07510_ (
    .A( dbg_0.dbg_reg_din_7_ ),
    .Y(_01025_)
  );
  INVX1 _07511_ (
    .A( dbg_0.dbg_reg_din_8_ ),
    .Y(_01026_)
  );
  INVX1 _07512_ (
    .A( dbg_0.dbg_reg_din_9_ ),
    .Y(_01027_)
  );
  INVX1 _07513_ (
    .A( dbg_0.dbg_reg_din_10_ ),
    .Y(_01028_)
  );
  INVX1 _07514_ (
    .A( dbg_0.dbg_reg_din_11_ ),
    .Y(_01029_)
  );
  INVX1 _07515_ (
    .A( dbg_0.dbg_reg_din_12_ ),
    .Y(_01030_)
  );
  INVX1 _07516_ (
    .A( dbg_0.dbg_reg_din_13_ ),
    .Y(_01031_)
  );
  INVX1 _07517_ (
    .A( dbg_0.dbg_reg_din_14_ ),
    .Y(_01032_)
  );
  INVX1 _07518_ (
    .A( dbg_0.dbg_reg_din_15_ ),
    .Y(_01033_)
  );
  INVX1 _07519_ (
    .A( execution_unit_0.inst_ad_6_ ),
    .Y(_01034_)
  );
  INVX1 _07520_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_01035_)
  );
  INVX1 _07521_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .Y(_01036_)
  );
  INVX1 _07522_ (
    .A( dbg_0.dbg_reg_wr ),
    .Y(_01037_)
  );
  INVX1 _07523_ (
    .A(_06327_),
    .Y(_00927_)
  );
  NOR2X1 _07524_ (
    .A( execution_unit_0.e_state_2_ ),
    .B(_01015_),
    .Y(_01038_)
  );
  AND2X1 _07525_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_01013_),
    .Y(_01039_)
  );
  NAND2X1 _07526_ (
    .A(_01038_),
    .B(_01039_),
    .Y(_01040_)
  );
  NOR2X1 _07527_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01040_),
    .Y(_01041_)
  );
  NAND3X1 _07528_ (
    .A(_01016_),
    .B(_01038_),
    .C(_01039_),
    .Y(_01042_)
  );
  AND2X1 _07529_ (
    .A( execution_unit_0.e_state_1_ ),
    .B( execution_unit_0.e_state_0_ ),
    .Y(_01043_)
  );
  NOR2X1 _07530_ (
    .A(_01014_),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_01044_)
  );
  NAND2X1 _07531_ (
    .A(_01043_),
    .B(_01044_),
    .Y(_01045_)
  );
  NOR2X1 _07532_ (
    .A( execution_unit_0.e_state_2_ ),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_01046_)
  );
  NAND2X1 _07533_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_01046_),
    .Y(_01047_)
  );
  OAI21X1 _07534_ (
    .A( execution_unit_0.inst_irq_rst ),
    .B(_01047_),
    .C(_01045_),
    .Y(_01048_)
  );
  OAI21X1 _07535_ (
    .A(_01041_),
    .B(_01048_),
    .C(_01036_),
    .Y(_01049_)
  );
  NAND3X1 _07536_ (
    .A( execution_unit_0.e_state_1_ ),
    .B( execution_unit_0.e_state_2_ ),
    .C(_01015_),
    .Y(_01050_)
  );
  OR2X1 _07537_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_01050_),
    .Y(_01051_)
  );
  INVX1 _07538_ (
    .A(_01051_),
    .Y(_00926_)
  );
  NOR2X1 _07539_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_01013_),
    .Y(_01052_)
  );
  AND2X1 _07540_ (
    .A(_01038_),
    .B(_01052_),
    .Y(_01053_)
  );
  NAND2X1 _07541_ (
    .A(_01038_),
    .B(_01052_),
    .Y(_01054_)
  );
  NOR2X1 _07542_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B( execution_unit_0.inst_mov ),
    .Y(_01055_)
  );
  NAND3X1 _07543_ (
    .A(_01014_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_01043_),
    .Y(_01056_)
  );
  INVX1 _07544_ (
    .A(_01056_),
    .Y( execution_unit_0.alu_0.exec_cycle )
  );
  NAND2X1 _07545_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01057_)
  );
  AOI22X1 _07546_ (
    .A(_01017_),
    .B(_00926_),
    .C(_01053_),
    .D(_01055_),
    .Y(_01058_)
  );
  NAND3X1 _07547_ (
    .A(_01049_),
    .B(_01057_),
    .C(_01058_),
    .Y( dbg_0.UNUSED_eu_mb_en )
  );
  MUX2X1 _07548_ (
    .A( dbg_0.UNUSED_eu_mab_0_ ),
    .B( execution_unit_0.mab_lsb ),
    .S( dbg_0.UNUSED_eu_mb_en ),
    .Y(_01059_)
  );
  INVX1 _07549_ (
    .A(_01059_),
    .Y(_00995_)
  );
  OAI21X1 _07550_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_en ),
    .C(_01056_),
    .Y(_01060_)
  );
  INVX1 _07551_ (
    .A(_01060_),
    .Y(_00994_)
  );
  NAND2X1 _07552_ (
    .A( execution_unit_0.mdb_in_15_ ),
    .B( execution_unit_0.mdb_in_buf_en ),
    .Y(_01061_)
  );
  OAI21X1 _07553_ (
    .A(_00997_),
    .B( execution_unit_0.mdb_in_buf_en ),
    .C(_01061_),
    .Y(_00993_)
  );
  NAND2X1 _07554_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_14_ ),
    .Y(_01062_)
  );
  OAI21X1 _07555_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00998_),
    .C(_01062_),
    .Y(_00992_)
  );
  NAND2X1 _07556_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_13_ ),
    .Y(_01063_)
  );
  OAI21X1 _07557_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00999_),
    .C(_01063_),
    .Y(_00991_)
  );
  NAND2X1 _07558_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_12_ ),
    .Y(_01064_)
  );
  OAI21X1 _07559_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01000_),
    .C(_01064_),
    .Y(_00990_)
  );
  NAND2X1 _07560_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_11_ ),
    .Y(_01065_)
  );
  OAI21X1 _07561_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01001_),
    .C(_01065_),
    .Y(_00989_)
  );
  NAND2X1 _07562_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_10_ ),
    .Y(_01066_)
  );
  OAI21X1 _07563_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01002_),
    .C(_01066_),
    .Y(_00988_)
  );
  NAND2X1 _07564_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_9_ ),
    .Y(_01067_)
  );
  OAI21X1 _07565_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01003_),
    .C(_01067_),
    .Y(_00987_)
  );
  NAND2X1 _07566_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_8_ ),
    .Y(_01068_)
  );
  OAI21X1 _07567_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01004_),
    .C(_01068_),
    .Y(_00986_)
  );
  NAND2X1 _07568_ (
    .A( execution_unit_0.mab_lsb ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01069_)
  );
  MUX2X1 _07569_ (
    .A( execution_unit_0.mdb_in_7_ ),
    .B( execution_unit_0.mdb_in_15_ ),
    .S(_01069_),
    .Y(_01070_)
  );
  NOR2X1 _07570_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_7_ ),
    .Y(_01071_)
  );
  AOI21X1 _07571_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01070_),
    .C(_01071_),
    .Y(_00985_)
  );
  MUX2X1 _07572_ (
    .A( execution_unit_0.mdb_in_6_ ),
    .B( execution_unit_0.mdb_in_14_ ),
    .S(_01069_),
    .Y(_01072_)
  );
  NOR2X1 _07573_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_6_ ),
    .Y(_01073_)
  );
  AOI21X1 _07574_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01072_),
    .C(_01073_),
    .Y(_00984_)
  );
  MUX2X1 _07575_ (
    .A( execution_unit_0.mdb_in_5_ ),
    .B( execution_unit_0.mdb_in_13_ ),
    .S(_01069_),
    .Y(_01074_)
  );
  NOR2X1 _07576_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_5_ ),
    .Y(_01075_)
  );
  AOI21X1 _07577_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01074_),
    .C(_01075_),
    .Y(_00983_)
  );
  MUX2X1 _07578_ (
    .A( execution_unit_0.mdb_in_4_ ),
    .B( execution_unit_0.mdb_in_12_ ),
    .S(_01069_),
    .Y(_01076_)
  );
  NOR2X1 _07579_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_4_ ),
    .Y(_01077_)
  );
  AOI21X1 _07580_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01076_),
    .C(_01077_),
    .Y(_00982_)
  );
  MUX2X1 _07581_ (
    .A( execution_unit_0.mdb_in_3_ ),
    .B( execution_unit_0.mdb_in_11_ ),
    .S(_01069_),
    .Y(_01078_)
  );
  NOR2X1 _07582_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_3_ ),
    .Y(_01079_)
  );
  AOI21X1 _07583_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01078_),
    .C(_01079_),
    .Y(_00981_)
  );
  MUX2X1 _07584_ (
    .A( execution_unit_0.mdb_in_2_ ),
    .B( execution_unit_0.mdb_in_10_ ),
    .S(_01069_),
    .Y(_01080_)
  );
  NOR2X1 _07585_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_2_ ),
    .Y(_01081_)
  );
  AOI21X1 _07586_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01080_),
    .C(_01081_),
    .Y(_00980_)
  );
  MUX2X1 _07587_ (
    .A( execution_unit_0.mdb_in_1_ ),
    .B( execution_unit_0.mdb_in_9_ ),
    .S(_01069_),
    .Y(_01082_)
  );
  NOR2X1 _07588_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_1_ ),
    .Y(_01083_)
  );
  AOI21X1 _07589_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01082_),
    .C(_01083_),
    .Y(_00979_)
  );
  MUX2X1 _07590_ (
    .A( execution_unit_0.mdb_in_0_ ),
    .B( execution_unit_0.mdb_in_8_ ),
    .S(_01069_),
    .Y(_01084_)
  );
  NOR2X1 _07591_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_0_ ),
    .Y(_01085_)
  );
  AOI21X1 _07592_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01084_),
    .C(_01085_),
    .Y(_00978_)
  );
  NAND2X1 _07593_ (
    .A(_01013_),
    .B(_01046_),
    .Y(_01086_)
  );
  OAI21X1 _07594_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_01056_),
    .C(_01054_),
    .Y(_01087_)
  );
  AOI21X1 _07595_ (
    .A(_01013_),
    .B(_01046_),
    .C(_01087_),
    .Y(_01088_)
  );
  MUX2X1 _07596_ (
    .A( execution_unit_0.pc_nxt_15_ ),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .S(_01053_),
    .Y(_01089_)
  );
  NAND2X1 _07597_ (
    .A( execution_unit_0.mdb_out_nxt_15_ ),
    .B(_01088_),
    .Y(_01090_)
  );
  OAI21X1 _07598_ (
    .A(_01088_),
    .B(_01089_),
    .C(_01090_),
    .Y(_00977_)
  );
  MUX2X1 _07599_ (
    .A( execution_unit_0.pc_nxt_14_ ),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .S(_01053_),
    .Y(_01091_)
  );
  NAND2X1 _07600_ (
    .A( execution_unit_0.mdb_out_nxt_14_ ),
    .B(_01088_),
    .Y(_01092_)
  );
  OAI21X1 _07601_ (
    .A(_01088_),
    .B(_01091_),
    .C(_01092_),
    .Y(_00976_)
  );
  MUX2X1 _07602_ (
    .A( execution_unit_0.pc_nxt_13_ ),
    .B( execution_unit_0.alu_0.alu_out_13_ ),
    .S(_01053_),
    .Y(_01093_)
  );
  NAND2X1 _07603_ (
    .A( execution_unit_0.mdb_out_nxt_13_ ),
    .B(_01088_),
    .Y(_01094_)
  );
  OAI21X1 _07604_ (
    .A(_01088_),
    .B(_01093_),
    .C(_01094_),
    .Y(_00975_)
  );
  MUX2X1 _07605_ (
    .A( execution_unit_0.pc_nxt_12_ ),
    .B( execution_unit_0.alu_0.alu_out_12_ ),
    .S(_01053_),
    .Y(_01095_)
  );
  NAND2X1 _07606_ (
    .A( execution_unit_0.mdb_out_nxt_12_ ),
    .B(_01088_),
    .Y(_01096_)
  );
  OAI21X1 _07607_ (
    .A(_01088_),
    .B(_01095_),
    .C(_01096_),
    .Y(_00974_)
  );
  MUX2X1 _07608_ (
    .A( execution_unit_0.pc_nxt_11_ ),
    .B( execution_unit_0.alu_0.alu_out_11_ ),
    .S(_01053_),
    .Y(_01097_)
  );
  NAND2X1 _07609_ (
    .A( execution_unit_0.mdb_out_nxt_11_ ),
    .B(_01088_),
    .Y(_01098_)
  );
  OAI21X1 _07610_ (
    .A(_01088_),
    .B(_01097_),
    .C(_01098_),
    .Y(_00973_)
  );
  MUX2X1 _07611_ (
    .A( execution_unit_0.pc_nxt_10_ ),
    .B( execution_unit_0.alu_0.alu_out_10_ ),
    .S(_01053_),
    .Y(_01099_)
  );
  NAND2X1 _07612_ (
    .A( execution_unit_0.mdb_out_nxt_10_ ),
    .B(_01088_),
    .Y(_01100_)
  );
  OAI21X1 _07613_ (
    .A(_01088_),
    .B(_01099_),
    .C(_01100_),
    .Y(_00972_)
  );
  MUX2X1 _07614_ (
    .A( execution_unit_0.pc_nxt_9_ ),
    .B( execution_unit_0.alu_0.alu_out_9_ ),
    .S(_01053_),
    .Y(_01101_)
  );
  NAND2X1 _07615_ (
    .A( execution_unit_0.mdb_out_nxt_9_ ),
    .B(_01088_),
    .Y(_01102_)
  );
  OAI21X1 _07616_ (
    .A(_01088_),
    .B(_01101_),
    .C(_01102_),
    .Y(_00971_)
  );
  MUX2X1 _07617_ (
    .A( execution_unit_0.pc_nxt_8_ ),
    .B( execution_unit_0.alu_0.alu_out_8_ ),
    .S(_01053_),
    .Y(_01103_)
  );
  NAND2X1 _07618_ (
    .A( execution_unit_0.mdb_out_nxt_8_ ),
    .B(_01088_),
    .Y(_01104_)
  );
  OAI21X1 _07619_ (
    .A(_01088_),
    .B(_01103_),
    .C(_01104_),
    .Y(_00970_)
  );
  MUX2X1 _07620_ (
    .A( execution_unit_0.pc_nxt_7_ ),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .S(_01053_),
    .Y(_01105_)
  );
  NAND2X1 _07621_ (
    .A( execution_unit_0.mdb_out_7_ ),
    .B(_01088_),
    .Y(_01106_)
  );
  OAI21X1 _07622_ (
    .A(_01088_),
    .B(_01105_),
    .C(_01106_),
    .Y(_00969_)
  );
  MUX2X1 _07623_ (
    .A( execution_unit_0.pc_nxt_6_ ),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .S(_01053_),
    .Y(_01107_)
  );
  NAND2X1 _07624_ (
    .A( execution_unit_0.mdb_out_6_ ),
    .B(_01088_),
    .Y(_01108_)
  );
  OAI21X1 _07625_ (
    .A(_01088_),
    .B(_01107_),
    .C(_01108_),
    .Y(_00968_)
  );
  MUX2X1 _07626_ (
    .A( execution_unit_0.pc_nxt_5_ ),
    .B( execution_unit_0.alu_0.alu_out_5_ ),
    .S(_01053_),
    .Y(_01109_)
  );
  NAND2X1 _07627_ (
    .A( execution_unit_0.mdb_out_5_ ),
    .B(_01088_),
    .Y(_01110_)
  );
  OAI21X1 _07628_ (
    .A(_01088_),
    .B(_01109_),
    .C(_01110_),
    .Y(_00967_)
  );
  MUX2X1 _07629_ (
    .A( execution_unit_0.pc_nxt_4_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .S(_01053_),
    .Y(_01111_)
  );
  NAND2X1 _07630_ (
    .A( execution_unit_0.mdb_out_4_ ),
    .B(_01088_),
    .Y(_01112_)
  );
  OAI21X1 _07631_ (
    .A(_01088_),
    .B(_01111_),
    .C(_01112_),
    .Y(_00966_)
  );
  MUX2X1 _07632_ (
    .A( execution_unit_0.pc_nxt_3_ ),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .S(_01053_),
    .Y(_01113_)
  );
  NAND2X1 _07633_ (
    .A( execution_unit_0.mdb_out_3_ ),
    .B(_01088_),
    .Y(_01114_)
  );
  OAI21X1 _07634_ (
    .A(_01088_),
    .B(_01113_),
    .C(_01114_),
    .Y(_00965_)
  );
  MUX2X1 _07635_ (
    .A( execution_unit_0.pc_nxt_2_ ),
    .B( execution_unit_0.alu_0.alu_out_2_ ),
    .S(_01053_),
    .Y(_01115_)
  );
  NAND2X1 _07636_ (
    .A( execution_unit_0.mdb_out_2_ ),
    .B(_01088_),
    .Y(_01116_)
  );
  OAI21X1 _07637_ (
    .A(_01088_),
    .B(_01115_),
    .C(_01116_),
    .Y(_00964_)
  );
  MUX2X1 _07638_ (
    .A( execution_unit_0.pc_nxt_1_ ),
    .B( execution_unit_0.alu_0.alu_out_1_ ),
    .S(_01053_),
    .Y(_01117_)
  );
  NAND2X1 _07639_ (
    .A( execution_unit_0.mdb_out_1_ ),
    .B(_01088_),
    .Y(_01118_)
  );
  OAI21X1 _07640_ (
    .A(_01088_),
    .B(_01117_),
    .C(_01118_),
    .Y(_00963_)
  );
  MUX2X1 _07641_ (
    .A( execution_unit_0.pc_nxt_0_ ),
    .B( execution_unit_0.alu_0.alu_out_0_ ),
    .S(_01053_),
    .Y(_01119_)
  );
  NAND2X1 _07642_ (
    .A( execution_unit_0.mdb_out_0_ ),
    .B(_01088_),
    .Y(_01120_)
  );
  OAI21X1 _07643_ (
    .A(_01088_),
    .B(_01119_),
    .C(_01120_),
    .Y(_00962_)
  );
  NOR2X1 _07644_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_01086_),
    .Y( execution_unit_0.reg_sr_clr )
  );
  NOR2X1 _07645_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_01056_),
    .Y(_01121_)
  );
  OAI21X1 _07646_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B(_01050_),
    .C(_01086_),
    .Y(_01122_)
  );
  AOI21X1 _07647_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B(_01121_),
    .C(_01122_),
    .Y(_01123_)
  );
  NOR2X1 _07648_ (
    .A( execution_unit_0.reg_src_0_ ),
    .B(_01123_),
    .Y(_01124_)
  );
  NOR2X1 _07649_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01125_)
  );
  OR2X1 _07650_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01126_)
  );
  NOR3X1 _07651_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_01013_),
    .C(_01125_),
    .Y(_01127_)
  );
  NOR2X1 _07652_ (
    .A(_01054_),
    .B(_01125_),
    .Y(_01128_)
  );
  NAND2X1 _07653_ (
    .A(_01038_),
    .B(_01127_),
    .Y(_01129_)
  );
  NAND3X1 _07654_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B(_01044_),
    .C(_01127_),
    .Y(_01130_)
  );
  AND2X1 _07655_ (
    .A(_01047_),
    .B(_01130_),
    .Y(_01131_)
  );
  AND2X1 _07656_ (
    .A(_01129_),
    .B(_01131_),
    .Y(_01132_)
  );
  NOR2X1 _07657_ (
    .A(_01016_),
    .B(_01054_),
    .Y( execution_unit_0.reg_sr_wr )
  );
  NOR2X1 _07658_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.inst_as_2_ ),
    .Y(_01133_)
  );
  OR2X1 _07659_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B( execution_unit_0.inst_as_1_ ),
    .Y(_01134_)
  );
  NOR2X1 _07660_ (
    .A( execution_unit_0.inst_as_4_ ),
    .B(_01134_),
    .Y(_01135_)
  );
  AOI21X1 _07661_ (
    .A(_01133_),
    .B(_01135_),
    .C(_01056_),
    .Y(_01136_)
  );
  NOR2X1 _07662_ (
    .A( execution_unit_0.reg_sr_wr ),
    .B(_01136_),
    .Y(_01137_)
  );
  AOI21X1 _07663_ (
    .A(_01042_),
    .B(_01054_),
    .C(_01126_),
    .Y(_01138_)
  );
  NOR2X1 _07664_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( execution_unit_0.inst_as_7_ ),
    .Y(_01139_)
  );
  NOR2X1 _07665_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B( execution_unit_0.inst_as_5_ ),
    .Y(_01140_)
  );
  AOI21X1 _07666_ (
    .A(_01139_),
    .B(_01140_),
    .C(_01056_),
    .Y(_01141_)
  );
  AOI22X1 _07667_ (
    .A( execution_unit_0.inst_dext_0_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_0_ ),
    .Y(_01142_)
  );
  NOR2X1 _07668_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01084_),
    .Y(_01143_)
  );
  AOI21X1 _07669_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_0_ ),
    .C(_01143_),
    .Y(_01144_)
  );
  MUX2X1 _07670_ (
    .A(_01142_),
    .B(_01144_),
    .S(_01137_),
    .Y(_01145_)
  );
  OAI21X1 _07671_ (
    .A(_01018_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01146_)
  );
  AOI21X1 _07672_ (
    .A(_01132_),
    .B(_01145_),
    .C(_01146_),
    .Y(_01147_)
  );
  NOR2X1 _07673_ (
    .A(_01124_),
    .B(_01147_),
    .Y( execution_unit_0.alu_0.alu_swpb_8_ )
  );
  NOR2X1 _07674_ (
    .A( execution_unit_0.reg_src_1_ ),
    .B(_01123_),
    .Y(_01148_)
  );
  AOI22X1 _07675_ (
    .A( execution_unit_0.inst_dext_1_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_1_ ),
    .Y(_01149_)
  );
  NOR2X1 _07676_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01082_),
    .Y(_01150_)
  );
  AOI21X1 _07677_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_1_ ),
    .C(_01150_),
    .Y(_01151_)
  );
  MUX2X1 _07678_ (
    .A(_01149_),
    .B(_01151_),
    .S(_01137_),
    .Y(_01152_)
  );
  OAI21X1 _07679_ (
    .A(_01019_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01153_)
  );
  AOI21X1 _07680_ (
    .A(_01132_),
    .B(_01152_),
    .C(_01153_),
    .Y(_01154_)
  );
  NOR2X1 _07681_ (
    .A(_01148_),
    .B(_01154_),
    .Y( execution_unit_0.alu_0.alu_shift_0_ )
  );
  NOR2X1 _07682_ (
    .A( execution_unit_0.reg_src_2_ ),
    .B(_01123_),
    .Y(_01155_)
  );
  AOI22X1 _07683_ (
    .A( execution_unit_0.inst_dext_2_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_2_ ),
    .Y(_01156_)
  );
  NOR2X1 _07684_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01080_),
    .Y(_01157_)
  );
  AOI21X1 _07685_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_2_ ),
    .C(_01157_),
    .Y(_01158_)
  );
  MUX2X1 _07686_ (
    .A(_01156_),
    .B(_01158_),
    .S(_01137_),
    .Y(_01159_)
  );
  OAI21X1 _07687_ (
    .A(_01020_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01160_)
  );
  AOI21X1 _07688_ (
    .A(_01132_),
    .B(_01159_),
    .C(_01160_),
    .Y(_01161_)
  );
  NOR2X1 _07689_ (
    .A(_01155_),
    .B(_01161_),
    .Y( execution_unit_0.alu_0.alu_shift_1_ )
  );
  NOR2X1 _07690_ (
    .A( execution_unit_0.reg_src_3_ ),
    .B(_01123_),
    .Y(_01162_)
  );
  AOI22X1 _07691_ (
    .A( execution_unit_0.inst_dext_3_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_3_ ),
    .Y(_01163_)
  );
  NOR2X1 _07692_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01078_),
    .Y(_01164_)
  );
  AOI21X1 _07693_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_3_ ),
    .C(_01164_),
    .Y(_01165_)
  );
  MUX2X1 _07694_ (
    .A(_01163_),
    .B(_01165_),
    .S(_01137_),
    .Y(_01166_)
  );
  OAI21X1 _07695_ (
    .A(_01021_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01167_)
  );
  AOI21X1 _07696_ (
    .A(_01132_),
    .B(_01166_),
    .C(_01167_),
    .Y(_01168_)
  );
  NOR2X1 _07697_ (
    .A(_01162_),
    .B(_01168_),
    .Y( execution_unit_0.alu_0.alu_shift_2_ )
  );
  NOR2X1 _07698_ (
    .A( execution_unit_0.reg_src_4_ ),
    .B(_01123_),
    .Y(_01169_)
  );
  AOI22X1 _07699_ (
    .A( execution_unit_0.inst_dext_4_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_4_ ),
    .Y(_01170_)
  );
  NOR2X1 _07700_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01076_),
    .Y(_01171_)
  );
  AOI21X1 _07701_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_4_ ),
    .C(_01171_),
    .Y(_01172_)
  );
  MUX2X1 _07702_ (
    .A(_01170_),
    .B(_01172_),
    .S(_01137_),
    .Y(_01173_)
  );
  OAI21X1 _07703_ (
    .A(_01022_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01174_)
  );
  AOI21X1 _07704_ (
    .A(_01132_),
    .B(_01173_),
    .C(_01174_),
    .Y(_01175_)
  );
  NOR2X1 _07705_ (
    .A(_01169_),
    .B(_01175_),
    .Y( execution_unit_0.alu_0.alu_shift_3_ )
  );
  NOR2X1 _07706_ (
    .A( execution_unit_0.reg_src_5_ ),
    .B(_01123_),
    .Y(_01176_)
  );
  AOI22X1 _07707_ (
    .A( execution_unit_0.inst_dext_5_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_5_ ),
    .Y(_01177_)
  );
  NOR2X1 _07708_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01074_),
    .Y(_01178_)
  );
  AOI21X1 _07709_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_5_ ),
    .C(_01178_),
    .Y(_01179_)
  );
  MUX2X1 _07710_ (
    .A(_01177_),
    .B(_01179_),
    .S(_01137_),
    .Y(_01180_)
  );
  OAI21X1 _07711_ (
    .A(_01023_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01181_)
  );
  AOI21X1 _07712_ (
    .A(_01132_),
    .B(_01180_),
    .C(_01181_),
    .Y(_01182_)
  );
  NOR2X1 _07713_ (
    .A(_01176_),
    .B(_01182_),
    .Y( execution_unit_0.alu_0.alu_shift_4_ )
  );
  NOR2X1 _07714_ (
    .A( execution_unit_0.reg_src_6_ ),
    .B(_01123_),
    .Y(_01183_)
  );
  AOI22X1 _07715_ (
    .A( execution_unit_0.inst_dext_6_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_6_ ),
    .Y(_01184_)
  );
  NOR2X1 _07716_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01072_),
    .Y(_01185_)
  );
  AOI21X1 _07717_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_6_ ),
    .C(_01185_),
    .Y(_01186_)
  );
  MUX2X1 _07718_ (
    .A(_01184_),
    .B(_01186_),
    .S(_01137_),
    .Y(_01187_)
  );
  OAI21X1 _07719_ (
    .A(_01024_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01188_)
  );
  AOI21X1 _07720_ (
    .A(_01132_),
    .B(_01187_),
    .C(_01188_),
    .Y(_01189_)
  );
  NOR2X1 _07721_ (
    .A(_01183_),
    .B(_01189_),
    .Y( execution_unit_0.alu_0.alu_shift_5_ )
  );
  NOR2X1 _07722_ (
    .A( execution_unit_0.reg_src_7_ ),
    .B(_01123_),
    .Y(_01190_)
  );
  AOI22X1 _07723_ (
    .A( execution_unit_0.inst_dext_7_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_7_ ),
    .Y(_01191_)
  );
  NOR2X1 _07724_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01070_),
    .Y(_01192_)
  );
  AOI21X1 _07725_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_7_ ),
    .C(_01192_),
    .Y(_01193_)
  );
  MUX2X1 _07726_ (
    .A(_01191_),
    .B(_01193_),
    .S(_01137_),
    .Y(_01194_)
  );
  OAI21X1 _07727_ (
    .A(_01025_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01195_)
  );
  AOI21X1 _07728_ (
    .A(_01132_),
    .B(_01194_),
    .C(_01195_),
    .Y(_01196_)
  );
  NOR2X1 _07729_ (
    .A(_01190_),
    .B(_01196_),
    .Y( execution_unit_0.alu_0.alu_shift_6_ )
  );
  NOR2X1 _07730_ (
    .A( execution_unit_0.reg_src_8_ ),
    .B(_01123_),
    .Y(_01197_)
  );
  AOI22X1 _07731_ (
    .A( execution_unit_0.inst_dext_8_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_8_ ),
    .Y(_01198_)
  );
  MUX2X1 _07732_ (
    .A( execution_unit_0.mdb_in_buf_8_ ),
    .B( execution_unit_0.mdb_in_8_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01199_)
  );
  MUX2X1 _07733_ (
    .A(_01198_),
    .B(_01199_),
    .S(_01137_),
    .Y(_01200_)
  );
  OAI21X1 _07734_ (
    .A(_01026_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01201_)
  );
  AOI21X1 _07735_ (
    .A(_01132_),
    .B(_01200_),
    .C(_01201_),
    .Y(_01202_)
  );
  NOR2X1 _07736_ (
    .A(_01197_),
    .B(_01202_),
    .Y( execution_unit_0.alu_0.alu_swpb_0_ )
  );
  NOR2X1 _07737_ (
    .A( execution_unit_0.reg_src_9_ ),
    .B(_01123_),
    .Y(_01203_)
  );
  AOI22X1 _07738_ (
    .A( execution_unit_0.inst_dext_9_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_9_ ),
    .Y(_01204_)
  );
  MUX2X1 _07739_ (
    .A( execution_unit_0.mdb_in_buf_9_ ),
    .B( execution_unit_0.mdb_in_9_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01205_)
  );
  MUX2X1 _07740_ (
    .A(_01204_),
    .B(_01205_),
    .S(_01137_),
    .Y(_01206_)
  );
  OAI21X1 _07741_ (
    .A(_01027_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01207_)
  );
  AOI21X1 _07742_ (
    .A(_01132_),
    .B(_01206_),
    .C(_01207_),
    .Y(_01208_)
  );
  NOR2X1 _07743_ (
    .A(_01203_),
    .B(_01208_),
    .Y( execution_unit_0.alu_0.alu_shift_8_ )
  );
  NOR2X1 _07744_ (
    .A( execution_unit_0.reg_src_10_ ),
    .B(_01123_),
    .Y(_01209_)
  );
  AOI22X1 _07745_ (
    .A( execution_unit_0.inst_dext_10_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_10_ ),
    .Y(_01210_)
  );
  MUX2X1 _07746_ (
    .A( execution_unit_0.mdb_in_buf_10_ ),
    .B( execution_unit_0.mdb_in_10_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01211_)
  );
  MUX2X1 _07747_ (
    .A(_01210_),
    .B(_01211_),
    .S(_01137_),
    .Y(_01212_)
  );
  OAI21X1 _07748_ (
    .A(_01028_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01213_)
  );
  AOI21X1 _07749_ (
    .A(_01132_),
    .B(_01212_),
    .C(_01213_),
    .Y(_01214_)
  );
  NOR2X1 _07750_ (
    .A(_01209_),
    .B(_01214_),
    .Y( execution_unit_0.alu_0.alu_shift_9_ )
  );
  NOR2X1 _07751_ (
    .A( execution_unit_0.reg_src_11_ ),
    .B(_01123_),
    .Y(_01215_)
  );
  AOI22X1 _07752_ (
    .A( execution_unit_0.inst_dext_11_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_11_ ),
    .Y(_01216_)
  );
  MUX2X1 _07753_ (
    .A( execution_unit_0.mdb_in_buf_11_ ),
    .B( execution_unit_0.mdb_in_11_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01217_)
  );
  MUX2X1 _07754_ (
    .A(_01216_),
    .B(_01217_),
    .S(_01137_),
    .Y(_01218_)
  );
  OAI21X1 _07755_ (
    .A(_01029_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01219_)
  );
  AOI21X1 _07756_ (
    .A(_01132_),
    .B(_01218_),
    .C(_01219_),
    .Y(_01220_)
  );
  NOR2X1 _07757_ (
    .A(_01215_),
    .B(_01220_),
    .Y( execution_unit_0.alu_0.alu_shift_10_ )
  );
  NOR2X1 _07758_ (
    .A( execution_unit_0.reg_src_12_ ),
    .B(_01123_),
    .Y(_01221_)
  );
  AOI22X1 _07759_ (
    .A( execution_unit_0.inst_dext_12_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_12_ ),
    .Y(_01222_)
  );
  MUX2X1 _07760_ (
    .A( execution_unit_0.mdb_in_buf_12_ ),
    .B( execution_unit_0.mdb_in_12_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01223_)
  );
  MUX2X1 _07761_ (
    .A(_01222_),
    .B(_01223_),
    .S(_01137_),
    .Y(_01224_)
  );
  OAI21X1 _07762_ (
    .A(_01030_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01225_)
  );
  AOI21X1 _07763_ (
    .A(_01132_),
    .B(_01224_),
    .C(_01225_),
    .Y(_01226_)
  );
  NOR2X1 _07764_ (
    .A(_01221_),
    .B(_01226_),
    .Y( execution_unit_0.alu_0.alu_shift_11_ )
  );
  NOR2X1 _07765_ (
    .A( execution_unit_0.reg_src_13_ ),
    .B(_01123_),
    .Y(_01227_)
  );
  AOI22X1 _07766_ (
    .A( execution_unit_0.inst_dext_13_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_13_ ),
    .Y(_01228_)
  );
  MUX2X1 _07767_ (
    .A( execution_unit_0.mdb_in_buf_13_ ),
    .B( execution_unit_0.mdb_in_13_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01229_)
  );
  MUX2X1 _07768_ (
    .A(_01228_),
    .B(_01229_),
    .S(_01137_),
    .Y(_01230_)
  );
  OAI21X1 _07769_ (
    .A(_01031_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01231_)
  );
  AOI21X1 _07770_ (
    .A(_01132_),
    .B(_01230_),
    .C(_01231_),
    .Y(_01232_)
  );
  NOR2X1 _07771_ (
    .A(_01227_),
    .B(_01232_),
    .Y( execution_unit_0.alu_0.alu_shift_12_ )
  );
  NOR2X1 _07772_ (
    .A( execution_unit_0.reg_src_14_ ),
    .B(_01123_),
    .Y(_01233_)
  );
  AOI22X1 _07773_ (
    .A( execution_unit_0.inst_dext_14_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_14_ ),
    .Y(_01234_)
  );
  MUX2X1 _07774_ (
    .A( execution_unit_0.mdb_in_buf_14_ ),
    .B( execution_unit_0.mdb_in_14_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01235_)
  );
  MUX2X1 _07775_ (
    .A(_01234_),
    .B(_01235_),
    .S(_01137_),
    .Y(_01236_)
  );
  OAI21X1 _07776_ (
    .A(_01032_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01237_)
  );
  AOI21X1 _07777_ (
    .A(_01132_),
    .B(_01236_),
    .C(_01237_),
    .Y(_01238_)
  );
  NOR2X1 _07778_ (
    .A(_01233_),
    .B(_01238_),
    .Y( execution_unit_0.alu_0.alu_shift_13_ )
  );
  NOR2X1 _07779_ (
    .A( execution_unit_0.reg_src_15_ ),
    .B(_01123_),
    .Y(_01239_)
  );
  AOI22X1 _07780_ (
    .A( execution_unit_0.inst_dext_15_ ),
    .B(_01138_),
    .C(_01141_),
    .D( execution_unit_0.inst_sext_15_ ),
    .Y(_01240_)
  );
  MUX2X1 _07781_ (
    .A( execution_unit_0.mdb_in_buf_15_ ),
    .B( execution_unit_0.mdb_in_15_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01241_)
  );
  MUX2X1 _07782_ (
    .A(_01240_),
    .B(_01241_),
    .S(_01137_),
    .Y(_01242_)
  );
  OAI21X1 _07783_ (
    .A(_01033_),
    .B(_01132_),
    .C(_01123_),
    .Y(_01243_)
  );
  AOI21X1 _07784_ (
    .A(_01132_),
    .B(_01242_),
    .C(_01243_),
    .Y(_01244_)
  );
  NOR2X1 _07785_ (
    .A(_01239_),
    .B(_01244_),
    .Y( execution_unit_0.alu_0.alu_shift_14_ )
  );
  OR2X1 _07786_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( execution_unit_0.inst_ad_0_ ),
    .Y(_01245_)
  );
  NOR2X1 _07787_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B(_01245_),
    .Y(_01246_)
  );
  INVX1 _07788_ (
    .A(_01246_),
    .Y(_01247_)
  );
  OR2X1 _07789_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01056_),
    .Y(_01248_)
  );
  NOR2X1 _07790_ (
    .A(_01246_),
    .B(_01248_),
    .Y(_01249_)
  );
  NOR2X1 _07791_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01126_),
    .Y(_01250_)
  );
  INVX1 _07792_ (
    .A(_01250_),
    .Y(_01251_)
  );
  OAI21X1 _07793_ (
    .A(_01054_),
    .B(_01251_),
    .C(_01040_),
    .Y(_01252_)
  );
  AOI21X1 _07794_ (
    .A(_01034_),
    .B(_01252_),
    .C(_01249_),
    .Y(_01253_)
  );
  NOR2X1 _07795_ (
    .A(_01247_),
    .B(_01248_),
    .Y(_01254_)
  );
  NOR2X1 _07796_ (
    .A(_01016_),
    .B(_01040_),
    .Y(_01255_)
  );
  NOR2X1 _07797_ (
    .A(_01254_),
    .B(_01255_),
    .Y(_01256_)
  );
  OAI22X1 _07798_ (
    .A(_01016_),
    .B(_01040_),
    .C(_01247_),
    .D(_01248_),
    .Y(_01257_)
  );
  NOR2X1 _07799_ (
    .A(_01253_),
    .B(_01257_),
    .Y(_01258_)
  );
  NOR2X1 _07800_ (
    .A(_01050_),
    .B(_01135_),
    .Y(_01259_)
  );
  OR2X1 _07801_ (
    .A(_01050_),
    .B(_01135_),
    .Y(_01260_)
  );
  NAND2X1 _07802_ (
    .A( execution_unit_0.inst_sext_0_ ),
    .B(_01259_),
    .Y(_01261_)
  );
  OAI21X1 _07803_ (
    .A(_01084_),
    .B(_01256_),
    .C(_01261_),
    .Y(_01262_)
  );
  AOI21X1 _07804_ (
    .A( dbg_0.dbg_reg_din_0_ ),
    .B(_01258_),
    .C(_01262_),
    .Y(_01263_)
  );
  NAND2X1 _07805_ (
    .A(_06309_),
    .B( dbg_0.cpu_stat_full_0_ ),
    .Y(_01264_)
  );
  OAI21X1 _07806_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01263_),
    .C(_01264_),
    .Y( execution_unit_0.alu_0.op_dst_0_ )
  );
  NAND2X1 _07807_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06316_),
    .Y(_01265_)
  );
  OAI21X1 _07808_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.inst_as_2_ ),
    .C( execution_unit_0.inst_src_1_ ),
    .Y(_01266_)
  );
  OR2X1 _07809_ (
    .A(_01125_),
    .B(_01266_),
    .Y(_01267_)
  );
  OAI21X1 _07810_ (
    .A(_01051_),
    .B(_01267_),
    .C(_01130_),
    .Y(_01268_)
  );
  OAI21X1 _07811_ (
    .A( execution_unit_0.e_state_1_ ),
    .B( execution_unit_0.e_state_0_ ),
    .C(_01046_),
    .Y(_01269_)
  );
  OAI21X1 _07812_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01129_),
    .C(_01269_),
    .Y(_01270_)
  );
  NOR3X1 _07813_ (
    .A(_01257_),
    .B(_01268_),
    .C(_01270_),
    .Y(_01271_)
  );
  OAI21X1 _07814_ (
    .A(_01019_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01272_)
  );
  OAI21X1 _07815_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01082_),
    .Y(_01273_)
  );
  AOI21X1 _07816_ (
    .A(_01272_),
    .B(_01273_),
    .C(_01259_),
    .Y(_01274_)
  );
  OAI21X1 _07817_ (
    .A( execution_unit_0.inst_sext_1_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01275_)
  );
  OAI21X1 _07818_ (
    .A(_01274_),
    .B(_01275_),
    .C(_01265_),
    .Y( execution_unit_0.alu_0.op_dst_1_ )
  );
  NAND2X1 _07819_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06317_),
    .Y(_01276_)
  );
  OAI21X1 _07820_ (
    .A(_01020_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01277_)
  );
  OAI21X1 _07821_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01080_),
    .Y(_01278_)
  );
  AOI21X1 _07822_ (
    .A(_01277_),
    .B(_01278_),
    .C(_01259_),
    .Y(_01279_)
  );
  OAI21X1 _07823_ (
    .A( execution_unit_0.inst_sext_2_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01280_)
  );
  OAI21X1 _07824_ (
    .A(_01279_),
    .B(_01280_),
    .C(_01276_),
    .Y( execution_unit_0.alu_0.op_dst_2_ )
  );
  NAND2X1 _07825_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06318_),
    .Y(_01281_)
  );
  OAI21X1 _07826_ (
    .A(_01021_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01282_)
  );
  OAI21X1 _07827_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01078_),
    .Y(_01283_)
  );
  AOI21X1 _07828_ (
    .A(_01282_),
    .B(_01283_),
    .C(_01259_),
    .Y(_01284_)
  );
  OAI21X1 _07829_ (
    .A( execution_unit_0.inst_sext_3_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01285_)
  );
  OAI21X1 _07830_ (
    .A(_01284_),
    .B(_01285_),
    .C(_01281_),
    .Y( execution_unit_0.alu_0.op_dst_3_ )
  );
  NAND2X1 _07831_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06319_),
    .Y(_01286_)
  );
  OAI21X1 _07832_ (
    .A(_01022_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01287_)
  );
  OAI21X1 _07833_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01076_),
    .Y(_01288_)
  );
  AOI21X1 _07834_ (
    .A(_01287_),
    .B(_01288_),
    .C(_01259_),
    .Y(_01289_)
  );
  OAI21X1 _07835_ (
    .A( execution_unit_0.inst_sext_4_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01290_)
  );
  OAI21X1 _07836_ (
    .A(_01289_),
    .B(_01290_),
    .C(_01286_),
    .Y( execution_unit_0.alu_0.op_dst_4_ )
  );
  NAND2X1 _07837_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06320_),
    .Y(_01291_)
  );
  OAI21X1 _07838_ (
    .A(_01023_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01292_)
  );
  OAI21X1 _07839_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01074_),
    .Y(_01293_)
  );
  AOI21X1 _07840_ (
    .A(_01292_),
    .B(_01293_),
    .C(_01259_),
    .Y(_01294_)
  );
  OAI21X1 _07841_ (
    .A( execution_unit_0.inst_sext_5_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01295_)
  );
  OAI21X1 _07842_ (
    .A(_01294_),
    .B(_01295_),
    .C(_01291_),
    .Y( execution_unit_0.alu_0.op_dst_5_ )
  );
  NAND2X1 _07843_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06321_),
    .Y(_01296_)
  );
  OAI21X1 _07844_ (
    .A(_01024_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01297_)
  );
  OAI21X1 _07845_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01072_),
    .Y(_01298_)
  );
  AOI21X1 _07846_ (
    .A(_01297_),
    .B(_01298_),
    .C(_01259_),
    .Y(_01299_)
  );
  OAI21X1 _07847_ (
    .A( execution_unit_0.inst_sext_6_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01300_)
  );
  OAI21X1 _07848_ (
    .A(_01299_),
    .B(_01300_),
    .C(_01296_),
    .Y( execution_unit_0.alu_0.op_dst_6_ )
  );
  NAND2X1 _07849_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06322_),
    .Y(_01301_)
  );
  OAI21X1 _07850_ (
    .A(_01025_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01302_)
  );
  OAI21X1 _07851_ (
    .A(_01254_),
    .B(_01255_),
    .C(_01070_),
    .Y(_01303_)
  );
  AOI21X1 _07852_ (
    .A(_01302_),
    .B(_01303_),
    .C(_01259_),
    .Y(_01304_)
  );
  OAI21X1 _07853_ (
    .A( execution_unit_0.inst_sext_7_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01305_)
  );
  OAI21X1 _07854_ (
    .A(_01304_),
    .B(_01305_),
    .C(_01301_),
    .Y( execution_unit_0.alu_0.op_dst_7_ )
  );
  NAND2X1 _07855_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06323_),
    .Y(_01306_)
  );
  OAI21X1 _07856_ (
    .A(_01026_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01307_)
  );
  OR2X1 _07857_ (
    .A( execution_unit_0.mdb_in_8_ ),
    .B(_01256_),
    .Y(_01308_)
  );
  AOI21X1 _07858_ (
    .A(_01307_),
    .B(_01308_),
    .C(_01259_),
    .Y(_01309_)
  );
  OAI21X1 _07859_ (
    .A( execution_unit_0.inst_sext_8_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01310_)
  );
  OAI21X1 _07860_ (
    .A(_01309_),
    .B(_01310_),
    .C(_01306_),
    .Y( execution_unit_0.alu_0.op_dst_8_ )
  );
  NAND2X1 _07861_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06324_),
    .Y(_01311_)
  );
  OAI21X1 _07862_ (
    .A(_01027_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01312_)
  );
  OR2X1 _07863_ (
    .A( execution_unit_0.mdb_in_9_ ),
    .B(_01256_),
    .Y(_01313_)
  );
  AOI21X1 _07864_ (
    .A(_01312_),
    .B(_01313_),
    .C(_01259_),
    .Y(_01314_)
  );
  OAI21X1 _07865_ (
    .A( execution_unit_0.inst_sext_9_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01315_)
  );
  OAI21X1 _07866_ (
    .A(_01314_),
    .B(_01315_),
    .C(_01311_),
    .Y( execution_unit_0.alu_0.op_dst_9_ )
  );
  NAND2X1 _07867_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06310_),
    .Y(_01316_)
  );
  OAI21X1 _07868_ (
    .A(_01028_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01317_)
  );
  OR2X1 _07869_ (
    .A( execution_unit_0.mdb_in_10_ ),
    .B(_01256_),
    .Y(_01318_)
  );
  AOI21X1 _07870_ (
    .A(_01317_),
    .B(_01318_),
    .C(_01259_),
    .Y(_01319_)
  );
  OAI21X1 _07871_ (
    .A( execution_unit_0.inst_sext_10_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01320_)
  );
  OAI21X1 _07872_ (
    .A(_01319_),
    .B(_01320_),
    .C(_01316_),
    .Y( execution_unit_0.alu_0.op_dst_10_ )
  );
  NAND2X1 _07873_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06311_),
    .Y(_01321_)
  );
  OAI21X1 _07874_ (
    .A(_01029_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01322_)
  );
  OR2X1 _07875_ (
    .A( execution_unit_0.mdb_in_11_ ),
    .B(_01256_),
    .Y(_01323_)
  );
  AOI21X1 _07876_ (
    .A(_01322_),
    .B(_01323_),
    .C(_01259_),
    .Y(_01324_)
  );
  OAI21X1 _07877_ (
    .A( execution_unit_0.inst_sext_11_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01325_)
  );
  OAI21X1 _07878_ (
    .A(_01324_),
    .B(_01325_),
    .C(_01321_),
    .Y( execution_unit_0.alu_0.op_dst_11_ )
  );
  NAND2X1 _07879_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06312_),
    .Y(_01326_)
  );
  OAI21X1 _07880_ (
    .A(_01030_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01327_)
  );
  OR2X1 _07881_ (
    .A( execution_unit_0.mdb_in_12_ ),
    .B(_01256_),
    .Y(_01328_)
  );
  AOI21X1 _07882_ (
    .A(_01327_),
    .B(_01328_),
    .C(_01259_),
    .Y(_01329_)
  );
  OAI21X1 _07883_ (
    .A( execution_unit_0.inst_sext_12_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01330_)
  );
  OAI21X1 _07884_ (
    .A(_01329_),
    .B(_01330_),
    .C(_01326_),
    .Y( execution_unit_0.alu_0.op_dst_12_ )
  );
  NAND2X1 _07885_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06313_),
    .Y(_01331_)
  );
  OAI21X1 _07886_ (
    .A(_01031_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01332_)
  );
  OR2X1 _07887_ (
    .A( execution_unit_0.mdb_in_13_ ),
    .B(_01256_),
    .Y(_01333_)
  );
  AOI21X1 _07888_ (
    .A(_01332_),
    .B(_01333_),
    .C(_01259_),
    .Y(_01334_)
  );
  OAI21X1 _07889_ (
    .A( execution_unit_0.inst_sext_13_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01335_)
  );
  OAI21X1 _07890_ (
    .A(_01334_),
    .B(_01335_),
    .C(_01331_),
    .Y( execution_unit_0.alu_0.op_dst_13_ )
  );
  NAND2X1 _07891_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06314_),
    .Y(_01336_)
  );
  OAI21X1 _07892_ (
    .A(_01032_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01337_)
  );
  OR2X1 _07893_ (
    .A( execution_unit_0.mdb_in_14_ ),
    .B(_01256_),
    .Y(_01338_)
  );
  AOI21X1 _07894_ (
    .A(_01337_),
    .B(_01338_),
    .C(_01259_),
    .Y(_01339_)
  );
  OAI21X1 _07895_ (
    .A( execution_unit_0.inst_sext_14_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01340_)
  );
  OAI21X1 _07896_ (
    .A(_01339_),
    .B(_01340_),
    .C(_01336_),
    .Y( execution_unit_0.alu_0.op_dst_14_ )
  );
  NAND2X1 _07897_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_06315_),
    .Y(_01341_)
  );
  OAI21X1 _07898_ (
    .A(_01033_),
    .B(_01253_),
    .C(_01271_),
    .Y(_01342_)
  );
  OR2X1 _07899_ (
    .A( execution_unit_0.mdb_in_15_ ),
    .B(_01256_),
    .Y(_01343_)
  );
  AOI21X1 _07900_ (
    .A(_01342_),
    .B(_01343_),
    .C(_01259_),
    .Y(_01344_)
  );
  OAI21X1 _07901_ (
    .A( execution_unit_0.inst_sext_15_ ),
    .B(_01260_),
    .C(_01035_),
    .Y(_01345_)
  );
  OAI21X1 _07902_ (
    .A(_01344_),
    .B(_01345_),
    .C(_01341_),
    .Y( execution_unit_0.alu_0.op_dst_15_ )
  );
  NAND2X1 _07903_ (
    .A( execution_unit_0.mdb_out_0_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01346_)
  );
  OAI21X1 _07904_ (
    .A(_01012_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01346_),
    .Y( execution_unit_0.mdb_out_8_ )
  );
  NAND2X1 _07905_ (
    .A( execution_unit_0.mdb_out_1_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01347_)
  );
  OAI21X1 _07906_ (
    .A(_01011_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01347_),
    .Y( execution_unit_0.mdb_out_9_ )
  );
  NAND2X1 _07907_ (
    .A( execution_unit_0.mdb_out_2_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01348_)
  );
  OAI21X1 _07908_ (
    .A(_01010_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01348_),
    .Y( execution_unit_0.mdb_out_10_ )
  );
  NAND2X1 _07909_ (
    .A( execution_unit_0.mdb_out_3_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01349_)
  );
  OAI21X1 _07910_ (
    .A(_01009_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01349_),
    .Y( execution_unit_0.mdb_out_11_ )
  );
  NAND2X1 _07911_ (
    .A( execution_unit_0.mdb_out_4_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01350_)
  );
  OAI21X1 _07912_ (
    .A(_01008_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01350_),
    .Y( execution_unit_0.mdb_out_12_ )
  );
  NAND2X1 _07913_ (
    .A( execution_unit_0.mdb_out_5_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01351_)
  );
  OAI21X1 _07914_ (
    .A(_01007_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01351_),
    .Y( execution_unit_0.mdb_out_13_ )
  );
  NAND2X1 _07915_ (
    .A( execution_unit_0.mdb_out_6_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01352_)
  );
  OAI21X1 _07916_ (
    .A(_01006_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01352_),
    .Y( execution_unit_0.mdb_out_14_ )
  );
  NAND2X1 _07917_ (
    .A( execution_unit_0.mdb_out_7_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01353_)
  );
  OAI21X1 _07918_ (
    .A(_01005_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01353_),
    .Y( execution_unit_0.mdb_out_15_ )
  );
  NAND3X1 _07919_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B( execution_unit_0.inst_type_0_ ),
    .C(_01250_),
    .Y(_01354_)
  );
  NAND2X1 _07920_ (
    .A( execution_unit_0.inst_ad_0_ ),
    .B( execution_unit_0.inst_type_2_ ),
    .Y(_01355_)
  );
  OAI21X1 _07921_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_01355_),
    .C(_01354_),
    .Y(_01356_)
  );
  OAI21X1 _07922_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_01356_),
    .C( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01357_)
  );
  NAND2X1 _07923_ (
    .A(_01037_),
    .B(_01357_),
    .Y( execution_unit_0.reg_dest_wr )
  );
  NAND2X1 _07924_ (
    .A(_01128_),
    .B(_01266_),
    .Y(_01358_)
  );
  NOR2X1 _07925_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B(_01358_),
    .Y(_01359_)
  );
  NOR2X1 _07926_ (
    .A(_01268_),
    .B(_01359_),
    .Y(_01360_)
  );
  OAI21X1 _07927_ (
    .A( execution_unit_0.inst_irq_rst ),
    .B(_01047_),
    .C(_01360_),
    .Y( execution_unit_0.reg_sp_wr )
  );
  NAND2X1 _07928_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01361_)
  );
  OAI21X1 _07929_ (
    .A(_01016_),
    .B(_01040_),
    .C(_01361_),
    .Y( execution_unit_0.reg_pc_call )
  );
  AOI22X1 _07930_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.exec_done ),
    .C( execution_unit_0.alu_0.exec_cycle ),
    .D( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01362_)
  );
  OAI21X1 _07931_ (
    .A(_01016_),
    .B(_01051_),
    .C(_01362_),
    .Y( execution_unit_0.reg_incr )
  );
  AOI21X1 _07932_ (
    .A( dbg_0.UNUSED_eu_mab_0_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01049_),
    .Y( dbg_0.UNUSED_eu_mb_wr_0_ )
  );
  AOI21X1 _07933_ (
    .A(_00996_),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C(_01049_),
    .Y( dbg_0.UNUSED_eu_mb_wr_1_ )
  );
  INVX1 _07934_ (
    .A(_06327_),
    .Y(_00928_)
  );
  INVX1 _07935_ (
    .A(_06327_),
    .Y(_00929_)
  );
  INVX1 _07936_ (
    .A(_06327_),
    .Y(_00930_)
  );
  INVX1 _07937_ (
    .A(_06327_),
    .Y(_00931_)
  );
  INVX1 _07938_ (
    .A(_06327_),
    .Y(_00932_)
  );
  INVX1 _07939_ (
    .A(_06327_),
    .Y(_00933_)
  );
  INVX1 _07940_ (
    .A(_06327_),
    .Y(_00934_)
  );
  INVX1 _07941_ (
    .A(_06327_),
    .Y(_00935_)
  );
  INVX1 _07942_ (
    .A(_06327_),
    .Y(_00936_)
  );
  INVX1 _07943_ (
    .A(_06327_),
    .Y(_00937_)
  );
  INVX1 _07944_ (
    .A(_06327_),
    .Y(_00938_)
  );
  INVX1 _07945_ (
    .A(_06327_),
    .Y(_00939_)
  );
  INVX1 _07946_ (
    .A(_06327_),
    .Y(_00940_)
  );
  INVX1 _07947_ (
    .A(_06327_),
    .Y(_00941_)
  );
  INVX1 _07948_ (
    .A(_06327_),
    .Y(_00942_)
  );
  INVX1 _07949_ (
    .A(_06327_),
    .Y(_00943_)
  );
  INVX1 _07950_ (
    .A(_06327_),
    .Y(_00944_)
  );
  INVX1 _07951_ (
    .A(_06327_),
    .Y(_00945_)
  );
  INVX1 _07952_ (
    .A(_06327_),
    .Y(_00946_)
  );
  INVX1 _07953_ (
    .A(_06327_),
    .Y(_00947_)
  );
  INVX1 _07954_ (
    .A(_06327_),
    .Y(_00948_)
  );
  INVX1 _07955_ (
    .A(_06327_),
    .Y(_00949_)
  );
  INVX1 _07956_ (
    .A(_06327_),
    .Y(_00950_)
  );
  INVX1 _07957_ (
    .A(_06327_),
    .Y(_00951_)
  );
  INVX1 _07958_ (
    .A(_06327_),
    .Y(_00952_)
  );
  INVX1 _07959_ (
    .A(_06327_),
    .Y(_00953_)
  );
  INVX1 _07960_ (
    .A(_06327_),
    .Y(_00954_)
  );
  INVX1 _07961_ (
    .A(_06327_),
    .Y(_00955_)
  );
  INVX1 _07962_ (
    .A(_06327_),
    .Y(_00956_)
  );
  INVX1 _07963_ (
    .A(_06327_),
    .Y(_00957_)
  );
  INVX1 _07964_ (
    .A(_06327_),
    .Y(_00958_)
  );
  INVX1 _07965_ (
    .A(_06327_),
    .Y(_00959_)
  );
  INVX1 _07966_ (
    .A(_06327_),
    .Y(_00960_)
  );
  INVX1 _07967_ (
    .A(_06327_),
    .Y(_00961_)
  );
  DFFSR _07968_ (
    .CLK(dco_clk),
    .D(_00962_),
    .Q( execution_unit_0.mdb_out_0_ ),
    .R(_00927_),
    .S(1'h1)
  );
  DFFSR _07969_ (
    .CLK(dco_clk),
    .D(_00963_),
    .Q( execution_unit_0.mdb_out_1_ ),
    .R(_00928_),
    .S(1'h1)
  );
  DFFSR _07970_ (
    .CLK(dco_clk),
    .D(_00964_),
    .Q( execution_unit_0.mdb_out_2_ ),
    .R(_00929_),
    .S(1'h1)
  );
  DFFSR _07971_ (
    .CLK(dco_clk),
    .D(_00965_),
    .Q( execution_unit_0.mdb_out_3_ ),
    .R(_00930_),
    .S(1'h1)
  );
  DFFSR _07972_ (
    .CLK(dco_clk),
    .D(_00966_),
    .Q( execution_unit_0.mdb_out_4_ ),
    .R(_00931_),
    .S(1'h1)
  );
  DFFSR _07973_ (
    .CLK(dco_clk),
    .D(_00967_),
    .Q( execution_unit_0.mdb_out_5_ ),
    .R(_00932_),
    .S(1'h1)
  );
  DFFSR _07974_ (
    .CLK(dco_clk),
    .D(_00968_),
    .Q( execution_unit_0.mdb_out_6_ ),
    .R(_00933_),
    .S(1'h1)
  );
  DFFSR _07975_ (
    .CLK(dco_clk),
    .D(_00969_),
    .Q( execution_unit_0.mdb_out_7_ ),
    .R(_00934_),
    .S(1'h1)
  );
  DFFSR _07976_ (
    .CLK(dco_clk),
    .D(_00970_),
    .Q( execution_unit_0.mdb_out_nxt_8_ ),
    .R(_00935_),
    .S(1'h1)
  );
  DFFSR _07977_ (
    .CLK(dco_clk),
    .D(_00971_),
    .Q( execution_unit_0.mdb_out_nxt_9_ ),
    .R(_00936_),
    .S(1'h1)
  );
  DFFSR _07978_ (
    .CLK(dco_clk),
    .D(_00972_),
    .Q( execution_unit_0.mdb_out_nxt_10_ ),
    .R(_00937_),
    .S(1'h1)
  );
  DFFSR _07979_ (
    .CLK(dco_clk),
    .D(_00973_),
    .Q( execution_unit_0.mdb_out_nxt_11_ ),
    .R(_00938_),
    .S(1'h1)
  );
  DFFSR _07980_ (
    .CLK(dco_clk),
    .D(_00974_),
    .Q( execution_unit_0.mdb_out_nxt_12_ ),
    .R(_00939_),
    .S(1'h1)
  );
  DFFSR _07981_ (
    .CLK(dco_clk),
    .D(_00975_),
    .Q( execution_unit_0.mdb_out_nxt_13_ ),
    .R(_00940_),
    .S(1'h1)
  );
  DFFSR _07982_ (
    .CLK(dco_clk),
    .D(_00976_),
    .Q( execution_unit_0.mdb_out_nxt_14_ ),
    .R(_00941_),
    .S(1'h1)
  );
  DFFSR _07983_ (
    .CLK(dco_clk),
    .D(_00977_),
    .Q( execution_unit_0.mdb_out_nxt_15_ ),
    .R(_00942_),
    .S(1'h1)
  );
  DFFSR _07984_ (
    .CLK(dco_clk),
    .D(_00978_),
    .Q( execution_unit_0.mdb_in_buf_0_ ),
    .R(_00943_),
    .S(1'h1)
  );
  DFFSR _07985_ (
    .CLK(dco_clk),
    .D(_00979_),
    .Q( execution_unit_0.mdb_in_buf_1_ ),
    .R(_00944_),
    .S(1'h1)
  );
  DFFSR _07986_ (
    .CLK(dco_clk),
    .D(_00980_),
    .Q( execution_unit_0.mdb_in_buf_2_ ),
    .R(_00945_),
    .S(1'h1)
  );
  DFFSR _07987_ (
    .CLK(dco_clk),
    .D(_00981_),
    .Q( execution_unit_0.mdb_in_buf_3_ ),
    .R(_00946_),
    .S(1'h1)
  );
  DFFSR _07988_ (
    .CLK(dco_clk),
    .D(_00982_),
    .Q( execution_unit_0.mdb_in_buf_4_ ),
    .R(_00947_),
    .S(1'h1)
  );
  DFFSR _07989_ (
    .CLK(dco_clk),
    .D(_00983_),
    .Q( execution_unit_0.mdb_in_buf_5_ ),
    .R(_00948_),
    .S(1'h1)
  );
  DFFSR _07990_ (
    .CLK(dco_clk),
    .D(_00984_),
    .Q( execution_unit_0.mdb_in_buf_6_ ),
    .R(_00949_),
    .S(1'h1)
  );
  DFFSR _07991_ (
    .CLK(dco_clk),
    .D(_00985_),
    .Q( execution_unit_0.mdb_in_buf_7_ ),
    .R(_00950_),
    .S(1'h1)
  );
  DFFSR _07992_ (
    .CLK(dco_clk),
    .D(_00986_),
    .Q( execution_unit_0.mdb_in_buf_8_ ),
    .R(_00951_),
    .S(1'h1)
  );
  DFFSR _07993_ (
    .CLK(dco_clk),
    .D(_00987_),
    .Q( execution_unit_0.mdb_in_buf_9_ ),
    .R(_00952_),
    .S(1'h1)
  );
  DFFSR _07994_ (
    .CLK(dco_clk),
    .D(_00988_),
    .Q( execution_unit_0.mdb_in_buf_10_ ),
    .R(_00953_),
    .S(1'h1)
  );
  DFFSR _07995_ (
    .CLK(dco_clk),
    .D(_00989_),
    .Q( execution_unit_0.mdb_in_buf_11_ ),
    .R(_00954_),
    .S(1'h1)
  );
  DFFSR _07996_ (
    .CLK(dco_clk),
    .D(_00990_),
    .Q( execution_unit_0.mdb_in_buf_12_ ),
    .R(_00955_),
    .S(1'h1)
  );
  DFFSR _07997_ (
    .CLK(dco_clk),
    .D(_00991_),
    .Q( execution_unit_0.mdb_in_buf_13_ ),
    .R(_00956_),
    .S(1'h1)
  );
  DFFSR _07998_ (
    .CLK(dco_clk),
    .D(_00992_),
    .Q( execution_unit_0.mdb_in_buf_14_ ),
    .R(_00957_),
    .S(1'h1)
  );
  DFFSR _07999_ (
    .CLK(dco_clk),
    .D(_00993_),
    .Q( execution_unit_0.mdb_in_buf_15_ ),
    .R(_00958_),
    .S(1'h1)
  );
  DFFSR _08000_ (
    .CLK(dco_clk),
    .D(_00926_),
    .Q( execution_unit_0.mdb_in_buf_en ),
    .R(_00959_),
    .S(1'h1)
  );
  DFFSR _08001_ (
    .CLK(dco_clk),
    .D(_00994_),
    .Q( execution_unit_0.mdb_in_buf_valid ),
    .R(_00960_),
    .S(1'h1)
  );
  DFFSR _08002_ (
    .CLK(dco_clk),
    .D(_00995_),
    .Q( execution_unit_0.mab_lsb ),
    .R(_00961_),
    .S(1'h1)
  );
  INVX1 _08003_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01899_)
  );
  INVX1 _08004_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01363_)
  );
  INVX1 _08005_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01364_)
  );
  INVX1 _08006_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01365_)
  );
  INVX1 _08007_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01366_)
  );
  INVX1 _08008_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .Y(_01367_)
  );
  INVX1 _08009_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01368_)
  );
  INVX1 _08010_ (
    .A( execution_unit_0.alu_0.inst_jmp_4_ ),
    .Y(_01369_)
  );
  INVX1 _08011_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .Y(_01370_)
  );
  INVX1 _08012_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .Y(_01371_)
  );
  OR2X1 _08013_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_01372_)
  );
  NOR2X1 _08014_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .Y(_01373_)
  );
  OR2X1 _08015_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .Y(_01374_)
  );
  AOI21X1 _08016_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.alu_0.inst_alu_2_ ),
    .C( execution_unit_0.alu_0.inst_alu_1_ ),
    .Y(_01375_)
  );
  NOR2X1 _08017_ (
    .A(_01899_),
    .B(_01375_),
    .Y(_01376_)
  );
  MUX2X1 _08018_ (
    .A( execution_unit_0.alu_0.inst_jmp_0_ ),
    .B( execution_unit_0.alu_0.inst_jmp_1_ ),
    .S( execution_unit_0.alu_0.status_1_ ),
    .Y(_01377_)
  );
  INVX1 _08019_ (
    .A(_01377_),
    .Y(_01378_)
  );
  MUX2X1 _08020_ (
    .A( execution_unit_0.alu_0.inst_jmp_2_ ),
    .B( execution_unit_0.alu_0.inst_jmp_3_ ),
    .S( execution_unit_0.alu_0.status_0_ ),
    .Y(_01379_)
  );
  OAI21X1 _08021_ (
    .A( execution_unit_0.alu_0.status_2_ ),
    .B(_01369_),
    .C(_01379_),
    .Y(_01380_)
  );
  NOR2X1 _08022_ (
    .A(_01378_),
    .B(_01380_),
    .Y(_01381_)
  );
  XOR2X1 _08023_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B( execution_unit_0.alu_0.status_2_ ),
    .Y(_01382_)
  );
  MUX2X1 _08024_ (
    .A( execution_unit_0.alu_0.inst_jmp_5_ ),
    .B( execution_unit_0.alu_0.inst_jmp_6_ ),
    .S(_01382_),
    .Y(_01383_)
  );
  AND2X1 _08025_ (
    .A(_01381_),
    .B(_01383_),
    .Y(_01384_)
  );
  NAND2X1 _08026_ (
    .A(_01381_),
    .B(_01383_),
    .Y(_01385_)
  );
  NAND2X1 _08027_ (
    .A( execution_unit_0.alu_0.inst_alu_0_ ),
    .B( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01386_)
  );
  XNOR2X1 _08028_ (
    .A( execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(_01386_),
    .Y(_01387_)
  );
  NOR2X1 _08029_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01387_),
    .Y(_01388_)
  );
  OR2X1 _08030_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01387_),
    .Y(_01389_)
  );
  AND2X1 _08031_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01387_),
    .Y(_01390_)
  );
  NAND2X1 _08032_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01387_),
    .Y(_01391_)
  );
  NAND2X1 _08033_ (
    .A(_01384_),
    .B(_01391_),
    .Y(_01392_)
  );
  OAI21X1 _08034_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01384_),
    .C(_01389_),
    .Y(_01393_)
  );
  AOI21X1 _08035_ (
    .A(_01384_),
    .B(_01390_),
    .C(_01393_),
    .Y( dbg_0.UNUSED_eu_mab_0_ )
  );
  NAND2X1 _08036_ (
    .A(_01376_),
    .B( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01394_)
  );
  XNOR2X1 _08037_ (
    .A(_01376_),
    .B( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01395_)
  );
  NAND2X1 _08038_ (
    .A(_01389_),
    .B(_01391_),
    .Y(_01396_)
  );
  OR2X1 _08039_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01397_)
  );
  NOR2X1 _08040_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01398_)
  );
  NAND3X1 _08041_ (
    .A(_01365_),
    .B(_01366_),
    .C(_01398_),
    .Y(_01399_)
  );
  NOR2X1 _08042_ (
    .A(_01397_),
    .B(_01399_),
    .Y(_01400_)
  );
  AOI21X1 _08043_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_swpb_0_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01401_)
  );
  AOI22X1 _08044_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_alu_10_ ),
    .C( execution_unit_0.alu_0.inst_so_3_ ),
    .D( execution_unit_0.alu_0.alu_swpb_8_ ),
    .Y(_01402_)
  );
  NAND2X1 _08045_ (
    .A(_01401_),
    .B(_01402_),
    .Y(_01403_)
  );
  AOI21X1 _08046_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01389_),
    .C(_01403_),
    .Y(_01404_)
  );
  AOI22X1 _08047_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01390_),
    .C(_01400_),
    .D(_01387_),
    .Y(_01405_)
  );
  AND2X1 _08048_ (
    .A(_01404_),
    .B(_01405_),
    .Y(_01406_)
  );
  OAI21X1 _08049_ (
    .A(_01365_),
    .B(_01396_),
    .C(_01406_),
    .Y(_01407_)
  );
  XNOR2X1 _08050_ (
    .A(_01367_),
    .B(_01396_),
    .Y(_01408_)
  );
  AOI21X1 _08051_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01408_),
    .C(_01374_),
    .Y(_01409_)
  );
  NAND2X1 _08052_ (
    .A(_01407_),
    .B(_01409_),
    .Y(_01410_)
  );
  OAI21X1 _08053_ (
    .A(_01373_),
    .B(_01395_),
    .C(_01410_),
    .Y( execution_unit_0.alu_0.alu_out_0_ )
  );
  XNOR2X1 _08054_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B(_01386_),
    .Y(_01411_)
  );
  NOR2X1 _08055_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01411_),
    .Y(_01412_)
  );
  AND2X1 _08056_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01411_),
    .Y(_01413_)
  );
  INVX1 _08057_ (
    .A(_01413_),
    .Y(_01414_)
  );
  NOR2X1 _08058_ (
    .A(_01412_),
    .B(_01413_),
    .Y(_01415_)
  );
  XNOR2X1 _08059_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01411_),
    .Y(_01416_)
  );
  NAND2X1 _08060_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01385_),
    .Y(_01417_)
  );
  NOR2X1 _08061_ (
    .A(_01391_),
    .B(_01416_),
    .Y(_01418_)
  );
  OAI21X1 _08062_ (
    .A(_01385_),
    .B(_01418_),
    .C(_01417_),
    .Y(_01419_)
  );
  OAI21X1 _08063_ (
    .A(_01392_),
    .B(_01415_),
    .C(_01419_),
    .Y(_01420_)
  );
  INVX1 _08064_ (
    .A(_01420_),
    .Y( dbg_0.UNUSED_eu_mab_1_ )
  );
  NOR2X1 _08065_ (
    .A(_01394_),
    .B(_01420_),
    .Y(_01421_)
  );
  NAND2X1 _08066_ (
    .A(_01394_),
    .B(_01420_),
    .Y(_01422_)
  );
  OAI21X1 _08067_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .C(_01422_),
    .Y(_01423_)
  );
  AOI21X1 _08068_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B(_01389_),
    .C(_01390_),
    .Y(_01424_)
  );
  OAI21X1 _08069_ (
    .A(_01367_),
    .B(_01388_),
    .C(_01391_),
    .Y(_01425_)
  );
  XNOR2X1 _08070_ (
    .A(_01415_),
    .B(_01424_),
    .Y(_01426_)
  );
  INVX1 _08071_ (
    .A(_01426_),
    .Y(_01427_)
  );
  XNOR2X1 _08072_ (
    .A( execution_unit_0.alu_0.alu_shift_2_ ),
    .B(_01386_),
    .Y(_01428_)
  );
  INVX1 _08073_ (
    .A(_01428_),
    .Y(_01429_)
  );
  NAND2X1 _08074_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01428_),
    .Y(_01430_)
  );
  INVX1 _08075_ (
    .A(_01430_),
    .Y(_01431_)
  );
  NAND2X1 _08076_ (
    .A(_01370_),
    .B(_01429_),
    .Y(_01432_)
  );
  NAND2X1 _08077_ (
    .A(_01430_),
    .B(_01432_),
    .Y(_01433_)
  );
  XNOR2X1 _08078_ (
    .A( execution_unit_0.alu_0.alu_shift_1_ ),
    .B(_01386_),
    .Y(_01434_)
  );
  AND2X1 _08079_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01434_),
    .Y(_01435_)
  );
  INVX1 _08080_ (
    .A(_01435_),
    .Y(_01436_)
  );
  AOI21X1 _08081_ (
    .A(_01415_),
    .B(_01425_),
    .C(_01413_),
    .Y(_01437_)
  );
  OAI21X1 _08082_ (
    .A(_01416_),
    .B(_01424_),
    .C(_01414_),
    .Y(_01438_)
  );
  NOR2X1 _08083_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01434_),
    .Y(_01439_)
  );
  INVX1 _08084_ (
    .A(_01439_),
    .Y(_01440_)
  );
  NAND2X1 _08085_ (
    .A(_01436_),
    .B(_01440_),
    .Y(_01441_)
  );
  AOI21X1 _08086_ (
    .A(_01438_),
    .B(_01440_),
    .C(_01435_),
    .Y(_01442_)
  );
  OAI21X1 _08087_ (
    .A(_01437_),
    .B(_01439_),
    .C(_01436_),
    .Y(_01443_)
  );
  AOI21X1 _08088_ (
    .A(_01432_),
    .B(_01443_),
    .C(_01431_),
    .Y(_01444_)
  );
  OAI21X1 _08089_ (
    .A(_01433_),
    .B(_01442_),
    .C(_01430_),
    .Y(_01445_)
  );
  XNOR2X1 _08090_ (
    .A(_01433_),
    .B(_01443_),
    .Y(_01446_)
  );
  XNOR2X1 _08091_ (
    .A(_01433_),
    .B(_01442_),
    .Y(_01447_)
  );
  XNOR2X1 _08092_ (
    .A(_01437_),
    .B(_01441_),
    .Y(_01448_)
  );
  AND2X1 _08093_ (
    .A(_01427_),
    .B(_01448_),
    .Y(_01449_)
  );
  NAND2X1 _08094_ (
    .A(_01427_),
    .B(_01448_),
    .Y(_01450_)
  );
  AOI21X1 _08095_ (
    .A(_01446_),
    .B(_01450_),
    .C(_01445_),
    .Y(_01451_)
  );
  OAI21X1 _08096_ (
    .A(_01447_),
    .B(_01449_),
    .C(_01444_),
    .Y(_01452_)
  );
  NOR2X1 _08097_ (
    .A(_01426_),
    .B(_01451_),
    .Y(_01453_)
  );
  OAI21X1 _08098_ (
    .A(_01427_),
    .B(_01452_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01454_)
  );
  OAI21X1 _08099_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01411_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01455_)
  );
  AOI22X1 _08100_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_1_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01456_)
  );
  NAND2X1 _08101_ (
    .A(_01368_),
    .B(_01456_),
    .Y(_01457_)
  );
  AOI21X1 _08102_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_8_ ),
    .C(_01457_),
    .Y(_01458_)
  );
  AOI22X1 _08103_ (
    .A(_01400_),
    .B(_01411_),
    .C(_01413_),
    .D( execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01459_)
  );
  NAND3X1 _08104_ (
    .A(_01455_),
    .B(_01458_),
    .C(_01459_),
    .Y(_01460_)
  );
  AOI21X1 _08105_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01415_),
    .C(_01460_),
    .Y(_01461_)
  );
  NOR2X1 _08106_ (
    .A(_01374_),
    .B(_01461_),
    .Y(_01462_)
  );
  OAI21X1 _08107_ (
    .A(_01453_),
    .B(_01454_),
    .C(_01462_),
    .Y(_01463_)
  );
  OAI21X1 _08108_ (
    .A(_01421_),
    .B(_01423_),
    .C(_01463_),
    .Y( execution_unit_0.alu_0.alu_out_1_ )
  );
  AOI21X1 _08109_ (
    .A(_01384_),
    .B(_01435_),
    .C(_01439_),
    .Y(_01464_)
  );
  OAI21X1 _08110_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01384_),
    .C(_01464_),
    .Y(_01465_)
  );
  OAI21X1 _08111_ (
    .A(_01413_),
    .B(_01418_),
    .C(_01384_),
    .Y(_01466_)
  );
  XOR2X1 _08112_ (
    .A(_01465_),
    .B(_01466_),
    .Y( dbg_0.UNUSED_eu_mab_2_ )
  );
  NAND2X1 _08113_ (
    .A(_01421_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_01467_)
  );
  XNOR2X1 _08114_ (
    .A(_01421_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_01468_)
  );
  NAND2X1 _08115_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01373_),
    .Y(_01469_)
  );
  NAND2X1 _08116_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_1_ ),
    .Y(_01470_)
  );
  AOI22X1 _08117_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C( execution_unit_0.alu_0.alu_shift_9_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01471_)
  );
  NAND3X1 _08118_ (
    .A(_01373_),
    .B(_01470_),
    .C(_01471_),
    .Y(_01472_)
  );
  AOI21X1 _08119_ (
    .A(_01400_),
    .B(_01434_),
    .C(_01472_),
    .Y(_01473_)
  );
  OAI21X1 _08120_ (
    .A(_01364_),
    .B(_01439_),
    .C(_01473_),
    .Y(_01474_)
  );
  AOI21X1 _08121_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01435_),
    .C(_01474_),
    .Y(_01475_)
  );
  OAI21X1 _08122_ (
    .A(_01365_),
    .B(_01441_),
    .C(_01475_),
    .Y(_01476_)
  );
  XNOR2X1 _08123_ (
    .A(_01448_),
    .B(_01453_),
    .Y(_01477_)
  );
  AOI22X1 _08124_ (
    .A(_01469_),
    .B(_01476_),
    .C(_01477_),
    .D( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01478_)
  );
  AOI21X1 _08125_ (
    .A(_01374_),
    .B(_01468_),
    .C(_01478_),
    .Y( execution_unit_0.alu_0.alu_out_2_ )
  );
  OAI22X1 _08126_ (
    .A(_01385_),
    .B(_01436_),
    .C(_01441_),
    .D(_01466_),
    .Y(_01479_)
  );
  OAI21X1 _08127_ (
    .A(_01385_),
    .B(_01429_),
    .C(_01370_),
    .Y(_01480_)
  );
  OAI21X1 _08128_ (
    .A(_01385_),
    .B(_01430_),
    .C(_01480_),
    .Y(_01481_)
  );
  XOR2X1 _08129_ (
    .A(_01479_),
    .B(_01481_),
    .Y(_01482_)
  );
  INVX1 _08130_ (
    .A(_01482_),
    .Y( dbg_0.UNUSED_eu_mab_3_ )
  );
  NOR2X1 _08131_ (
    .A(_01467_),
    .B(_01482_),
    .Y(_01483_)
  );
  XNOR2X1 _08132_ (
    .A(_01467_),
    .B(_01482_),
    .Y(_01484_)
  );
  OAI21X1 _08133_ (
    .A(_01444_),
    .B(_01449_),
    .C(_01447_),
    .Y(_01485_)
  );
  AND2X1 _08134_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01485_),
    .Y(_01486_)
  );
  OAI21X1 _08135_ (
    .A(_01447_),
    .B(_01449_),
    .C(_01486_),
    .Y(_01487_)
  );
  OAI21X1 _08136_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01428_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01488_)
  );
  AOI22X1 _08137_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C( execution_unit_0.alu_0.alu_shift_3_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01489_)
  );
  AOI22X1 _08138_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_10_ ),
    .C(_01400_),
    .D(_01428_),
    .Y(_01490_)
  );
  OAI21X1 _08139_ (
    .A(_01363_),
    .B(_01430_),
    .C(_01490_),
    .Y(_01491_)
  );
  INVX1 _08140_ (
    .A(_01491_),
    .Y(_01492_)
  );
  NAND3X1 _08141_ (
    .A(_01488_),
    .B(_01489_),
    .C(_01492_),
    .Y(_01493_)
  );
  OAI21X1 _08142_ (
    .A(_01365_),
    .B(_01433_),
    .C(_01373_),
    .Y(_01494_)
  );
  OAI21X1 _08143_ (
    .A(_01493_),
    .B(_01494_),
    .C(_01469_),
    .Y(_01495_)
  );
  AOI22X1 _08144_ (
    .A(_01374_),
    .B(_01484_),
    .C(_01487_),
    .D(_01495_),
    .Y( execution_unit_0.alu_0.alu_out_3_ )
  );
  XNOR2X1 _08145_ (
    .A( execution_unit_0.alu_0.alu_shift_3_ ),
    .B(_01386_),
    .Y(_01496_)
  );
  AND2X1 _08146_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01496_),
    .Y(_01497_)
  );
  NAND2X1 _08147_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01496_),
    .Y(_01498_)
  );
  NAND2X1 _08148_ (
    .A(_01384_),
    .B(_01496_),
    .Y(_01499_)
  );
  XOR2X1 _08149_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01499_),
    .Y(_01500_)
  );
  AOI22X1 _08150_ (
    .A(_01384_),
    .B(_01431_),
    .C(_01479_),
    .D(_01480_),
    .Y(_01501_)
  );
  XOR2X1 _08151_ (
    .A(_01500_),
    .B(_01501_),
    .Y( dbg_0.UNUSED_eu_mab_4_ )
  );
  NOR2X1 _08152_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01496_),
    .Y(_01502_)
  );
  NOR2X1 _08153_ (
    .A(_01497_),
    .B(_01502_),
    .Y(_01503_)
  );
  INVX1 _08154_ (
    .A(_01503_),
    .Y(_01504_)
  );
  NOR3X1 _08155_ (
    .A(_01444_),
    .B(_01447_),
    .C(_01449_),
    .Y(_01505_)
  );
  NAND3X1 _08156_ (
    .A(_01445_),
    .B(_01446_),
    .C(_01450_),
    .Y(_01506_)
  );
  OAI21X1 _08157_ (
    .A(_01451_),
    .B(_01505_),
    .C(_01504_),
    .Y(_01507_)
  );
  NOR3X1 _08158_ (
    .A(_01451_),
    .B(_01504_),
    .C(_01505_),
    .Y(_01508_)
  );
  NAND3X1 _08159_ (
    .A(_01452_),
    .B(_01503_),
    .C(_01506_),
    .Y(_01509_)
  );
  AND2X1 _08160_ (
    .A(_01507_),
    .B(_01509_),
    .Y(_01510_)
  );
  NAND2X1 _08161_ (
    .A(_01483_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_01511_)
  );
  XNOR2X1 _08162_ (
    .A(_01483_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_01512_)
  );
  AOI21X1 _08163_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_3_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01513_)
  );
  AOI22X1 _08164_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_11_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01514_)
  );
  NAND3X1 _08165_ (
    .A(_01373_),
    .B(_01513_),
    .C(_01514_),
    .Y(_01515_)
  );
  AOI21X1 _08166_ (
    .A(_01400_),
    .B(_01496_),
    .C(_01515_),
    .Y(_01516_)
  );
  OAI21X1 _08167_ (
    .A(_01364_),
    .B(_01502_),
    .C(_01516_),
    .Y(_01517_)
  );
  AOI21X1 _08168_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01497_),
    .C(_01517_),
    .Y(_01518_)
  );
  OAI21X1 _08169_ (
    .A(_01365_),
    .B(_01504_),
    .C(_01518_),
    .Y(_01519_)
  );
  OAI21X1 _08170_ (
    .A(_01469_),
    .B(_01510_),
    .C(_01519_),
    .Y(_01520_)
  );
  AOI21X1 _08171_ (
    .A(_01374_),
    .B(_01512_),
    .C(_01520_),
    .Y( execution_unit_0.alu_0.alu_out_4_ )
  );
  OAI22X1 _08172_ (
    .A(_01385_),
    .B(_01498_),
    .C(_01500_),
    .D(_01501_),
    .Y(_01521_)
  );
  INVX1 _08173_ (
    .A(_01521_),
    .Y(_01522_)
  );
  XNOR2X1 _08174_ (
    .A( execution_unit_0.alu_0.alu_shift_4_ ),
    .B(_01386_),
    .Y(_01523_)
  );
  AND2X1 _08175_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01523_),
    .Y(_01524_)
  );
  NAND2X1 _08176_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01523_),
    .Y(_01525_)
  );
  NOR2X1 _08177_ (
    .A(_01385_),
    .B(_01525_),
    .Y(_01526_)
  );
  AOI21X1 _08178_ (
    .A(_01384_),
    .B(_01523_),
    .C( execution_unit_0.alu_0.op_dst_5_ ),
    .Y(_01527_)
  );
  OR2X1 _08179_ (
    .A(_01526_),
    .B(_01527_),
    .Y(_01528_)
  );
  NOR2X1 _08180_ (
    .A(_01522_),
    .B(_01528_),
    .Y(_01529_)
  );
  XOR2X1 _08181_ (
    .A(_01521_),
    .B(_01528_),
    .Y(_01530_)
  );
  INVX1 _08182_ (
    .A(_01530_),
    .Y( dbg_0.UNUSED_eu_mab_5_ )
  );
  NOR2X1 _08183_ (
    .A(_01511_),
    .B(_01530_),
    .Y(_01531_)
  );
  INVX1 _08184_ (
    .A(_01531_),
    .Y(_01532_)
  );
  AOI21X1 _08185_ (
    .A(_01511_),
    .B(_01530_),
    .C(_01373_),
    .Y(_01533_)
  );
  OR2X1 _08186_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01523_),
    .Y(_01534_)
  );
  AND2X1 _08187_ (
    .A(_01525_),
    .B(_01534_),
    .Y(_01535_)
  );
  NAND2X1 _08188_ (
    .A(_01525_),
    .B(_01534_),
    .Y(_01536_)
  );
  AOI21X1 _08189_ (
    .A(_01498_),
    .B(_01509_),
    .C(_01536_),
    .Y(_01537_)
  );
  OAI21X1 _08190_ (
    .A(_01497_),
    .B(_01508_),
    .C(_01535_),
    .Y(_01538_)
  );
  NAND3X1 _08191_ (
    .A(_01498_),
    .B(_01509_),
    .C(_01536_),
    .Y(_01539_)
  );
  NAND2X1 _08192_ (
    .A(_01538_),
    .B(_01539_),
    .Y(_01540_)
  );
  XNOR2X1 _08193_ (
    .A( execution_unit_0.alu_0.alu_shift_5_ ),
    .B(_01386_),
    .Y(_01541_)
  );
  AND2X1 _08194_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01541_),
    .Y(_01542_)
  );
  NAND2X1 _08195_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01541_),
    .Y(_01543_)
  );
  XNOR2X1 _08196_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01541_),
    .Y(_01544_)
  );
  INVX1 _08197_ (
    .A(_01544_),
    .Y(_01545_)
  );
  NOR2X1 _08198_ (
    .A(_01524_),
    .B(_01537_),
    .Y(_01546_)
  );
  AOI21X1 _08199_ (
    .A(_01525_),
    .B(_01538_),
    .C(_01544_),
    .Y(_01547_)
  );
  OAI21X1 _08200_ (
    .A(_01524_),
    .B(_01537_),
    .C(_01545_),
    .Y(_01548_)
  );
  XNOR2X1 _08201_ (
    .A(_01544_),
    .B(_01546_),
    .Y(_01549_)
  );
  NAND2X1 _08202_ (
    .A(_01540_),
    .B(_01549_),
    .Y(_01550_)
  );
  OAI21X1 _08203_ (
    .A(_01544_),
    .B(_01546_),
    .C(_01543_),
    .Y(_01551_)
  );
  XNOR2X1 _08204_ (
    .A( execution_unit_0.alu_0.alu_shift_6_ ),
    .B(_01386_),
    .Y(_01552_)
  );
  AND2X1 _08205_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01552_),
    .Y(_01553_)
  );
  NAND2X1 _08206_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01552_),
    .Y(_01554_)
  );
  OR2X1 _08207_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01552_),
    .Y(_01555_)
  );
  NAND2X1 _08208_ (
    .A(_01554_),
    .B(_01555_),
    .Y(_01556_)
  );
  INVX1 _08209_ (
    .A(_01556_),
    .Y(_01557_)
  );
  NAND3X1 _08210_ (
    .A(_01543_),
    .B(_01548_),
    .C(_01557_),
    .Y(_01558_)
  );
  OAI21X1 _08211_ (
    .A(_01542_),
    .B(_01547_),
    .C(_01556_),
    .Y(_01559_)
  );
  NAND2X1 _08212_ (
    .A(_01558_),
    .B(_01559_),
    .Y(_01560_)
  );
  AOI22X1 _08213_ (
    .A(_01540_),
    .B(_01549_),
    .C(_01558_),
    .D(_01559_),
    .Y(_01561_)
  );
  NAND2X1 _08214_ (
    .A(_01550_),
    .B(_01560_),
    .Y(_01562_)
  );
  OAI21X1 _08215_ (
    .A(_01551_),
    .B(_01553_),
    .C(_01555_),
    .Y(_01563_)
  );
  NAND2X1 _08216_ (
    .A(_01562_),
    .B(_01563_),
    .Y(_01564_)
  );
  NAND2X1 _08217_ (
    .A(_01540_),
    .B(_01564_),
    .Y(_01565_)
  );
  XOR2X1 _08218_ (
    .A(_01540_),
    .B(_01564_),
    .Y(_01566_)
  );
  AOI21X1 _08219_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01567_)
  );
  AOI22X1 _08220_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_12_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01568_)
  );
  NAND2X1 _08221_ (
    .A(_01567_),
    .B(_01568_),
    .Y(_01569_)
  );
  AOI21X1 _08222_ (
    .A(_01400_),
    .B(_01523_),
    .C(_01569_),
    .Y(_01570_)
  );
  OAI21X1 _08223_ (
    .A(_01363_),
    .B(_01525_),
    .C(_01570_),
    .Y(_01571_)
  );
  AOI21X1 _08224_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01534_),
    .C(_01571_),
    .Y(_01572_)
  );
  OAI21X1 _08225_ (
    .A(_01365_),
    .B(_01536_),
    .C(_01572_),
    .Y(_01573_)
  );
  NAND2X1 _08226_ (
    .A(_01373_),
    .B(_01573_),
    .Y(_01574_)
  );
  AOI21X1 _08227_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01566_),
    .C(_01574_),
    .Y(_01575_)
  );
  AOI21X1 _08228_ (
    .A(_01532_),
    .B(_01533_),
    .C(_01575_),
    .Y(_01576_)
  );
  INVX1 _08229_ (
    .A(_01576_),
    .Y( execution_unit_0.alu_0.alu_out_5_ )
  );
  NOR2X1 _08230_ (
    .A(_01526_),
    .B(_01529_),
    .Y(_01577_)
  );
  NOR2X1 _08231_ (
    .A(_01385_),
    .B(_01543_),
    .Y(_01578_)
  );
  AOI21X1 _08232_ (
    .A(_01384_),
    .B(_01541_),
    .C( execution_unit_0.alu_0.op_dst_6_ ),
    .Y(_01579_)
  );
  OR2X1 _08233_ (
    .A(_01578_),
    .B(_01579_),
    .Y(_01580_)
  );
  OAI21X1 _08234_ (
    .A(_01578_),
    .B(_01579_),
    .C(_01577_),
    .Y(_01581_)
  );
  OR2X1 _08235_ (
    .A(_01577_),
    .B(_01580_),
    .Y(_01582_)
  );
  NAND2X1 _08236_ (
    .A(_01581_),
    .B(_01582_),
    .Y(_01583_)
  );
  INVX1 _08237_ (
    .A(_01583_),
    .Y( dbg_0.UNUSED_eu_mab_6_ )
  );
  NOR2X1 _08238_ (
    .A(_01532_),
    .B(_01583_),
    .Y(_01584_)
  );
  XOR2X1 _08239_ (
    .A(_01531_),
    .B(_01583_),
    .Y(_01585_)
  );
  OAI21X1 _08240_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01541_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01586_)
  );
  NAND2X1 _08241_ (
    .A(_01400_),
    .B(_01541_),
    .Y(_01587_)
  );
  AOI22X1 _08242_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C( execution_unit_0.alu_0.alu_shift_13_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01588_)
  );
  NAND2X1 _08243_ (
    .A(_01373_),
    .B(_01588_),
    .Y(_01589_)
  );
  AOI21X1 _08244_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C(_01589_),
    .Y(_01590_)
  );
  NAND2X1 _08245_ (
    .A(_01586_),
    .B(_01587_),
    .Y(_01591_)
  );
  OAI21X1 _08246_ (
    .A(_01365_),
    .B(_01544_),
    .C(_01590_),
    .Y(_01592_)
  );
  NOR2X1 _08247_ (
    .A(_01591_),
    .B(_01592_),
    .Y(_01593_)
  );
  OAI21X1 _08248_ (
    .A(_01363_),
    .B(_01543_),
    .C(_01593_),
    .Y(_01594_)
  );
  XOR2X1 _08249_ (
    .A(_01549_),
    .B(_01565_),
    .Y(_01595_)
  );
  AOI22X1 _08250_ (
    .A(_01469_),
    .B(_01594_),
    .C(_01595_),
    .D( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01596_)
  );
  AOI21X1 _08251_ (
    .A(_01374_),
    .B(_01585_),
    .C(_01596_),
    .Y( execution_unit_0.alu_0.alu_out_6_ )
  );
  AOI21X1 _08252_ (
    .A(_01550_),
    .B(_01555_),
    .C(_01560_),
    .Y(_01597_)
  );
  NOR2X1 _08253_ (
    .A(_01561_),
    .B(_01597_),
    .Y(_01598_)
  );
  OAI21X1 _08254_ (
    .A(_01385_),
    .B(_01543_),
    .C(_01582_),
    .Y(_01599_)
  );
  NOR2X1 _08255_ (
    .A(_01385_),
    .B(_01554_),
    .Y(_01600_)
  );
  OAI21X1 _08256_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01384_),
    .C(_01555_),
    .Y(_01601_)
  );
  NOR2X1 _08257_ (
    .A(_01600_),
    .B(_01601_),
    .Y(_01602_)
  );
  XOR2X1 _08258_ (
    .A(_01599_),
    .B(_01602_),
    .Y( dbg_0.UNUSED_eu_mab_7_ )
  );
  NAND2X1 _08259_ (
    .A(_01584_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01603_)
  );
  XNOR2X1 _08260_ (
    .A(_01584_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01604_)
  );
  OAI21X1 _08261_ (
    .A(_01365_),
    .B(_01553_),
    .C(_01364_),
    .Y(_01605_)
  );
  OAI21X1 _08262_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01552_),
    .C(_01605_),
    .Y(_01606_)
  );
  MUX2X1 _08263_ (
    .A( execution_unit_0.alu_0.alu_shift_6_ ),
    .B( execution_unit_0.alu_0.alu_shift_14_ ),
    .S( execution_unit_0.alu_0.inst_bw ),
    .Y(_01607_)
  );
  NOR2X1 _08264_ (
    .A( execution_unit_0.alu_0.inst_so_0_ ),
    .B(_01607_),
    .Y(_01608_)
  );
  AOI21X1 _08265_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.alu_0.inst_so_0_ ),
    .C(_01608_),
    .Y(_01609_)
  );
  OAI21X1 _08266_ (
    .A( execution_unit_0.alu_0.alu_swpb_0_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01610_)
  );
  AOI21X1 _08267_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01609_),
    .C(_01610_),
    .Y(_01611_)
  );
  AOI21X1 _08268_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01612_)
  );
  AOI21X1 _08269_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01374_),
    .Y(_01613_)
  );
  NAND2X1 _08270_ (
    .A(_01612_),
    .B(_01613_),
    .Y(_01614_)
  );
  AOI21X1 _08271_ (
    .A(_01400_),
    .B(_01552_),
    .C(_01614_),
    .Y(_01615_)
  );
  OAI21X1 _08272_ (
    .A(_01363_),
    .B(_01554_),
    .C(_01615_),
    .Y(_01616_)
  );
  NOR2X1 _08273_ (
    .A(_01611_),
    .B(_01616_),
    .Y(_01617_)
  );
  AOI22X1 _08274_ (
    .A(_01374_),
    .B(_01604_),
    .C(_01606_),
    .D(_01617_),
    .Y(_01618_)
  );
  OAI21X1 _08275_ (
    .A(_01469_),
    .B(_01598_),
    .C(_01618_),
    .Y(_01619_)
  );
  INVX1 _08276_ (
    .A(_01619_),
    .Y( execution_unit_0.alu_0.alu_out_7_ )
  );
  AOI21X1 _08277_ (
    .A(_01555_),
    .B(_01578_),
    .C(_01600_),
    .Y(_01620_)
  );
  OAI21X1 _08278_ (
    .A(_01582_),
    .B(_01601_),
    .C(_01620_),
    .Y(_01621_)
  );
  NOR2X1 _08279_ (
    .A(_01899_),
    .B(_01371_),
    .Y(_01622_)
  );
  NAND2X1 _08280_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01623_)
  );
  XOR2X1 _08281_ (
    .A( execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01386_),
    .Y(_01624_)
  );
  NOR2X1 _08282_ (
    .A(_01622_),
    .B(_01624_),
    .Y(_01625_)
  );
  OAI21X1 _08283_ (
    .A(_01899_),
    .B(_01371_),
    .C( execution_unit_0.alu_0.op_dst_8_ ),
    .Y(_01626_)
  );
  NOR2X1 _08284_ (
    .A(_01624_),
    .B(_01626_),
    .Y(_01627_)
  );
  INVX1 _08285_ (
    .A(_01627_),
    .Y(_01628_)
  );
  NAND2X1 _08286_ (
    .A(_01384_),
    .B(_01627_),
    .Y(_01629_)
  );
  AOI21X1 _08287_ (
    .A( execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01623_),
    .C(_01625_),
    .Y(_01630_)
  );
  AOI21X1 _08288_ (
    .A(_01385_),
    .B(_01626_),
    .C(_01630_),
    .Y(_01631_)
  );
  AND2X1 _08289_ (
    .A(_01629_),
    .B(_01631_),
    .Y(_01632_)
  );
  NAND2X1 _08290_ (
    .A(_01621_),
    .B(_01632_),
    .Y(_01633_)
  );
  XNOR2X1 _08291_ (
    .A(_01621_),
    .B(_01632_),
    .Y(_01634_)
  );
  INVX1 _08292_ (
    .A(_01634_),
    .Y( dbg_0.UNUSED_eu_mab_8_ )
  );
  NOR2X1 _08293_ (
    .A(_01627_),
    .B(_01630_),
    .Y(_01635_)
  );
  XNOR2X1 _08294_ (
    .A(_01561_),
    .B(_01563_),
    .Y(_01636_)
  );
  XOR2X1 _08295_ (
    .A(_01561_),
    .B(_01563_),
    .Y(_01637_)
  );
  XNOR2X1 _08296_ (
    .A(_01635_),
    .B(_01636_),
    .Y(_01638_)
  );
  AND2X1 _08297_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01635_),
    .Y(_01639_)
  );
  NAND2X1 _08298_ (
    .A(_01400_),
    .B(_01625_),
    .Y(_01640_)
  );
  AOI22X1 _08299_ (
    .A( execution_unit_0.alu_0.alu_swpb_8_ ),
    .B( execution_unit_0.alu_0.inst_so_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_8_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01641_)
  );
  NAND3X1 _08300_ (
    .A(_01612_),
    .B(_01640_),
    .C(_01641_),
    .Y(_01642_)
  );
  AOI21X1 _08301_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01627_),
    .C(_01642_),
    .Y(_01643_)
  );
  OAI21X1 _08302_ (
    .A(_01364_),
    .B(_01630_),
    .C(_01643_),
    .Y(_01644_)
  );
  OAI21X1 _08303_ (
    .A(_01639_),
    .B(_01644_),
    .C(_01373_),
    .Y(_01645_)
  );
  AOI21X1 _08304_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01638_),
    .C(_01645_),
    .Y(_01646_)
  );
  INVX1 _08305_ (
    .A(_01646_),
    .Y(_01647_)
  );
  AOI21X1 _08306_ (
    .A(_01584_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .C( dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_01648_)
  );
  OR2X1 _08307_ (
    .A(_01603_),
    .B(_01634_),
    .Y(_01649_)
  );
  OAI21X1 _08308_ (
    .A(_01603_),
    .B(_01634_),
    .C(_01374_),
    .Y(_01650_)
  );
  OAI21X1 _08309_ (
    .A(_01648_),
    .B(_01650_),
    .C(_01647_),
    .Y( execution_unit_0.alu_0.alu_out_8_ )
  );
  INVX1 _08310_ (
    .A( execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_01651_)
  );
  OAI21X1 _08311_ (
    .A(_01385_),
    .B(_01628_),
    .C(_01633_),
    .Y(_01652_)
  );
  XOR2X1 _08312_ (
    .A( execution_unit_0.alu_0.alu_shift_8_ ),
    .B(_01386_),
    .Y(_01653_)
  );
  NOR2X1 _08313_ (
    .A(_01622_),
    .B(_01653_),
    .Y(_01654_)
  );
  AND2X1 _08314_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01654_),
    .Y(_01655_)
  );
  NAND2X1 _08315_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01654_),
    .Y(_01656_)
  );
  NOR2X1 _08316_ (
    .A(_01385_),
    .B(_01656_),
    .Y(_01657_)
  );
  AOI21X1 _08317_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01623_),
    .C(_01654_),
    .Y(_01658_)
  );
  AOI22X1 _08318_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01623_),
    .C(_01654_),
    .D(_01384_),
    .Y(_01659_)
  );
  NOR2X1 _08319_ (
    .A(_01657_),
    .B(_01659_),
    .Y(_01660_)
  );
  XNOR2X1 _08320_ (
    .A(_01652_),
    .B(_01660_),
    .Y(_01661_)
  );
  INVX1 _08321_ (
    .A(_01661_),
    .Y( dbg_0.UNUSED_eu_mab_9_ )
  );
  AND2X1 _08322_ (
    .A(_01649_),
    .B(_01661_),
    .Y(_01662_)
  );
  OR2X1 _08323_ (
    .A(_01649_),
    .B(_01661_),
    .Y(_01663_)
  );
  OAI21X1 _08324_ (
    .A(_01649_),
    .B(_01661_),
    .C(_01374_),
    .Y(_01664_)
  );
  NOR2X1 _08325_ (
    .A(_01655_),
    .B(_01658_),
    .Y(_01665_)
  );
  AOI21X1 _08326_ (
    .A(_01635_),
    .B(_01636_),
    .C(_01627_),
    .Y(_01666_)
  );
  OAI21X1 _08327_ (
    .A(_01630_),
    .B(_01637_),
    .C(_01628_),
    .Y(_01667_)
  );
  XNOR2X1 _08328_ (
    .A(_01665_),
    .B(_01666_),
    .Y(_01668_)
  );
  XOR2X1 _08329_ (
    .A( execution_unit_0.alu_0.alu_shift_10_ ),
    .B(_01386_),
    .Y(_01669_)
  );
  NOR2X1 _08330_ (
    .A(_01622_),
    .B(_01669_),
    .Y(_01670_)
  );
  OAI21X1 _08331_ (
    .A(_01899_),
    .B(_01371_),
    .C( execution_unit_0.alu_0.op_dst_11_ ),
    .Y(_01671_)
  );
  NOR2X1 _08332_ (
    .A(_01669_),
    .B(_01671_),
    .Y(_01672_)
  );
  NAND2X1 _08333_ (
    .A( execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01670_),
    .Y(_01673_)
  );
  AOI21X1 _08334_ (
    .A( execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01623_),
    .C(_01670_),
    .Y(_01674_)
  );
  NOR2X1 _08335_ (
    .A(_01672_),
    .B(_01674_),
    .Y(_01675_)
  );
  XOR2X1 _08336_ (
    .A( execution_unit_0.alu_0.alu_shift_9_ ),
    .B(_01386_),
    .Y(_01676_)
  );
  NOR2X1 _08337_ (
    .A(_01622_),
    .B(_01676_),
    .Y(_01677_)
  );
  AND2X1 _08338_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01677_),
    .Y(_01678_)
  );
  INVX1 _08339_ (
    .A(_01678_),
    .Y(_01679_)
  );
  AOI21X1 _08340_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01623_),
    .C(_01677_),
    .Y(_01680_)
  );
  NOR2X1 _08341_ (
    .A(_01678_),
    .B(_01680_),
    .Y(_01681_)
  );
  AOI21X1 _08342_ (
    .A(_01665_),
    .B(_01667_),
    .C(_01655_),
    .Y(_01682_)
  );
  OAI21X1 _08343_ (
    .A(_01658_),
    .B(_01666_),
    .C(_01656_),
    .Y(_01683_)
  );
  AOI21X1 _08344_ (
    .A(_01681_),
    .B(_01683_),
    .C(_01678_),
    .Y(_01684_)
  );
  OAI21X1 _08345_ (
    .A(_01680_),
    .B(_01682_),
    .C(_01679_),
    .Y(_01685_)
  );
  AOI21X1 _08346_ (
    .A(_01675_),
    .B(_01685_),
    .C(_01672_),
    .Y(_01686_)
  );
  OAI21X1 _08347_ (
    .A(_01674_),
    .B(_01684_),
    .C(_01673_),
    .Y(_01687_)
  );
  XNOR2X1 _08348_ (
    .A(_01675_),
    .B(_01684_),
    .Y(_01688_)
  );
  XNOR2X1 _08349_ (
    .A(_01675_),
    .B(_01685_),
    .Y(_01689_)
  );
  XNOR2X1 _08350_ (
    .A(_01681_),
    .B(_01682_),
    .Y(_01690_)
  );
  NOR2X1 _08351_ (
    .A(_01668_),
    .B(_01690_),
    .Y(_01691_)
  );
  OR2X1 _08352_ (
    .A(_01668_),
    .B(_01690_),
    .Y(_01692_)
  );
  AOI21X1 _08353_ (
    .A(_01688_),
    .B(_01692_),
    .C(_01687_),
    .Y(_01693_)
  );
  OAI21X1 _08354_ (
    .A(_01689_),
    .B(_01691_),
    .C(_01686_),
    .Y(_01694_)
  );
  XNOR2X1 _08355_ (
    .A(_01668_),
    .B(_01693_),
    .Y(_01695_)
  );
  NAND2X1 _08356_ (
    .A(_01400_),
    .B(_01654_),
    .Y(_01696_)
  );
  AOI22X1 _08357_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_so_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_9_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01697_)
  );
  NAND3X1 _08358_ (
    .A(_01612_),
    .B(_01696_),
    .C(_01697_),
    .Y(_01698_)
  );
  AOI21X1 _08359_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01655_),
    .C(_01698_),
    .Y(_01699_)
  );
  OAI21X1 _08360_ (
    .A(_01364_),
    .B(_01658_),
    .C(_01699_),
    .Y(_01700_)
  );
  AOI21X1 _08361_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01665_),
    .C(_01700_),
    .Y(_01701_)
  );
  NOR2X1 _08362_ (
    .A(_01374_),
    .B(_01701_),
    .Y(_01702_)
  );
  OAI21X1 _08363_ (
    .A(_01368_),
    .B(_01695_),
    .C(_01702_),
    .Y(_01703_)
  );
  OAI21X1 _08364_ (
    .A(_01662_),
    .B(_01664_),
    .C(_01703_),
    .Y( execution_unit_0.alu_0.alu_out_9_ )
  );
  INVX1 _08365_ (
    .A( execution_unit_0.alu_0.alu_out_9_ ),
    .Y(_01704_)
  );
  NOR2X1 _08366_ (
    .A(_01629_),
    .B(_01658_),
    .Y(_01705_)
  );
  NOR2X1 _08367_ (
    .A(_01657_),
    .B(_01705_),
    .Y(_01706_)
  );
  OAI21X1 _08368_ (
    .A(_01633_),
    .B(_01659_),
    .C(_01706_),
    .Y(_01707_)
  );
  AOI22X1 _08369_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01623_),
    .C(_01677_),
    .D(_01384_),
    .Y(_01708_)
  );
  AOI21X1 _08370_ (
    .A(_01384_),
    .B(_01678_),
    .C(_01708_),
    .Y(_01709_)
  );
  NAND2X1 _08371_ (
    .A(_01707_),
    .B(_01709_),
    .Y(_01710_)
  );
  XNOR2X1 _08372_ (
    .A(_01707_),
    .B(_01709_),
    .Y(_01711_)
  );
  INVX1 _08373_ (
    .A(_01711_),
    .Y( dbg_0.UNUSED_eu_mab_10_ )
  );
  NOR2X1 _08374_ (
    .A(_01663_),
    .B(_01711_),
    .Y(_01712_)
  );
  OAI21X1 _08375_ (
    .A(_01649_),
    .B(_01661_),
    .C(_01711_),
    .Y(_01713_)
  );
  OAI21X1 _08376_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .C(_01713_),
    .Y(_01714_)
  );
  OAI21X1 _08377_ (
    .A(_01668_),
    .B(_01693_),
    .C(_01690_),
    .Y(_01715_)
  );
  AOI21X1 _08378_ (
    .A(_01687_),
    .B(_01691_),
    .C(_01368_),
    .Y(_01716_)
  );
  NAND2X1 _08379_ (
    .A(_01715_),
    .B(_01716_),
    .Y(_01717_)
  );
  NAND2X1 _08380_ (
    .A(_01400_),
    .B(_01677_),
    .Y(_01718_)
  );
  AOI22X1 _08381_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_10_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01719_)
  );
  NAND3X1 _08382_ (
    .A(_01612_),
    .B(_01718_),
    .C(_01719_),
    .Y(_01720_)
  );
  AOI21X1 _08383_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01678_),
    .C(_01720_),
    .Y(_01721_)
  );
  OAI21X1 _08384_ (
    .A(_01364_),
    .B(_01680_),
    .C(_01721_),
    .Y(_01722_)
  );
  AOI21X1 _08385_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01681_),
    .C(_01722_),
    .Y(_01723_)
  );
  NOR2X1 _08386_ (
    .A(_01374_),
    .B(_01723_),
    .Y(_01724_)
  );
  NAND2X1 _08387_ (
    .A(_01717_),
    .B(_01724_),
    .Y(_01725_)
  );
  OAI21X1 _08388_ (
    .A(_01712_),
    .B(_01714_),
    .C(_01725_),
    .Y( execution_unit_0.alu_0.alu_out_10_ )
  );
  NAND2X1 _08389_ (
    .A(_01384_),
    .B(_01670_),
    .Y(_01726_)
  );
  AOI22X1 _08390_ (
    .A(_01384_),
    .B(_01672_),
    .C(_01726_),
    .D(_01671_),
    .Y(_01727_)
  );
  OAI21X1 _08391_ (
    .A(_01385_),
    .B(_01679_),
    .C(_01710_),
    .Y(_01728_)
  );
  NAND2X1 _08392_ (
    .A(_01727_),
    .B(_01728_),
    .Y(_01729_)
  );
  XOR2X1 _08393_ (
    .A(_01727_),
    .B(_01728_),
    .Y( dbg_0.UNUSED_eu_mab_11_ )
  );
  NAND2X1 _08394_ (
    .A(_01712_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_01730_)
  );
  XOR2X1 _08395_ (
    .A(_01712_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_01731_)
  );
  AOI22X1 _08396_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_11_ ),
    .C( execution_unit_0.alu_0.alu_shift_6_ ),
    .D( execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01732_)
  );
  AOI22X1 _08397_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C(_01400_),
    .D(_01670_),
    .Y(_01733_)
  );
  OAI21X1 _08398_ (
    .A(_01363_),
    .B(_01673_),
    .C(_01733_),
    .Y(_01734_)
  );
  OAI21X1 _08399_ (
    .A(_01364_),
    .B(_01674_),
    .C(_01732_),
    .Y(_01735_)
  );
  NOR2X1 _08400_ (
    .A(_01734_),
    .B(_01735_),
    .Y(_01736_)
  );
  AOI21X1 _08401_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01675_),
    .C(_01374_),
    .Y(_01737_)
  );
  AOI22X1 _08402_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01373_),
    .C(_01736_),
    .D(_01737_),
    .Y(_01738_)
  );
  AOI21X1 _08403_ (
    .A(_01687_),
    .B(_01692_),
    .C(_01688_),
    .Y(_01739_)
  );
  OAI21X1 _08404_ (
    .A(_01689_),
    .B(_01691_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01740_)
  );
  NOR2X1 _08405_ (
    .A(_01739_),
    .B(_01740_),
    .Y(_01741_)
  );
  OAI22X1 _08406_ (
    .A(_01373_),
    .B(_01731_),
    .C(_01738_),
    .D(_01741_),
    .Y(_01742_)
  );
  INVX1 _08407_ (
    .A(_01742_),
    .Y( execution_unit_0.alu_0.alu_out_11_ )
  );
  OAI21X1 _08408_ (
    .A(_01385_),
    .B(_01673_),
    .C(_01729_),
    .Y(_01743_)
  );
  XOR2X1 _08409_ (
    .A( execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01386_),
    .Y(_01744_)
  );
  NOR2X1 _08410_ (
    .A(_01622_),
    .B(_01744_),
    .Y(_01745_)
  );
  AND2X1 _08411_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01745_),
    .Y(_01746_)
  );
  NAND2X1 _08412_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01745_),
    .Y(_01747_)
  );
  NAND2X1 _08413_ (
    .A(_01384_),
    .B(_01746_),
    .Y(_01748_)
  );
  AOI21X1 _08414_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01623_),
    .C(_01745_),
    .Y(_01749_)
  );
  AOI22X1 _08415_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01623_),
    .C(_01745_),
    .D(_01384_),
    .Y(_01750_)
  );
  AOI21X1 _08416_ (
    .A(_01384_),
    .B(_01746_),
    .C(_01750_),
    .Y(_01751_)
  );
  NAND2X1 _08417_ (
    .A(_01743_),
    .B(_01751_),
    .Y(_01752_)
  );
  XNOR2X1 _08418_ (
    .A(_01743_),
    .B(_01751_),
    .Y(_01753_)
  );
  INVX1 _08419_ (
    .A(_01753_),
    .Y( dbg_0.UNUSED_eu_mab_12_ )
  );
  NOR2X1 _08420_ (
    .A(_01730_),
    .B(_01753_),
    .Y(_01754_)
  );
  NAND2X1 _08421_ (
    .A(_01730_),
    .B(_01753_),
    .Y(_01755_)
  );
  OAI21X1 _08422_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .C(_01755_),
    .Y(_01756_)
  );
  NOR2X1 _08423_ (
    .A(_01746_),
    .B(_01749_),
    .Y(_01757_)
  );
  INVX1 _08424_ (
    .A(_01757_),
    .Y(_01758_)
  );
  NOR3X1 _08425_ (
    .A(_01686_),
    .B(_01689_),
    .C(_01691_),
    .Y(_01759_)
  );
  NAND3X1 _08426_ (
    .A(_01687_),
    .B(_01688_),
    .C(_01692_),
    .Y(_01760_)
  );
  OAI21X1 _08427_ (
    .A(_01693_),
    .B(_01759_),
    .C(_01758_),
    .Y(_01761_)
  );
  NOR3X1 _08428_ (
    .A(_01693_),
    .B(_01758_),
    .C(_01759_),
    .Y(_01762_)
  );
  NAND3X1 _08429_ (
    .A(_01694_),
    .B(_01757_),
    .C(_01760_),
    .Y(_01763_)
  );
  AND2X1 _08430_ (
    .A(_01761_),
    .B(_01763_),
    .Y(_01764_)
  );
  NAND2X1 _08431_ (
    .A(_01400_),
    .B(_01745_),
    .Y(_01765_)
  );
  AOI22X1 _08432_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_12_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01766_)
  );
  NAND3X1 _08433_ (
    .A(_01612_),
    .B(_01765_),
    .C(_01766_),
    .Y(_01767_)
  );
  AOI21X1 _08434_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01746_),
    .C(_01767_),
    .Y(_01768_)
  );
  OAI21X1 _08435_ (
    .A(_01364_),
    .B(_01749_),
    .C(_01768_),
    .Y(_01769_)
  );
  AOI21X1 _08436_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01757_),
    .C(_01769_),
    .Y(_01770_)
  );
  NOR2X1 _08437_ (
    .A(_01374_),
    .B(_01770_),
    .Y(_01771_)
  );
  OAI21X1 _08438_ (
    .A(_01368_),
    .B(_01764_),
    .C(_01771_),
    .Y(_01772_)
  );
  OAI21X1 _08439_ (
    .A(_01754_),
    .B(_01756_),
    .C(_01772_),
    .Y( execution_unit_0.alu_0.alu_out_12_ )
  );
  OAI21X1 _08440_ (
    .A(_01385_),
    .B(_01747_),
    .C(_01752_),
    .Y(_01773_)
  );
  XOR2X1 _08441_ (
    .A( execution_unit_0.alu_0.alu_shift_12_ ),
    .B(_01386_),
    .Y(_01774_)
  );
  NOR2X1 _08442_ (
    .A(_01622_),
    .B(_01774_),
    .Y(_01775_)
  );
  AND2X1 _08443_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01775_),
    .Y(_01776_)
  );
  NAND2X1 _08444_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01775_),
    .Y(_01777_)
  );
  AOI21X1 _08445_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01623_),
    .C(_01775_),
    .Y(_01778_)
  );
  AOI22X1 _08446_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01623_),
    .C(_01775_),
    .D(_01384_),
    .Y(_01779_)
  );
  AOI21X1 _08447_ (
    .A(_01384_),
    .B(_01776_),
    .C(_01779_),
    .Y(_01780_)
  );
  XOR2X1 _08448_ (
    .A(_01773_),
    .B(_01780_),
    .Y( dbg_0.UNUSED_eu_mab_13_ )
  );
  AND2X1 _08449_ (
    .A(_01754_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01781_)
  );
  XNOR2X1 _08450_ (
    .A(_01754_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01782_)
  );
  NOR2X1 _08451_ (
    .A(_01776_),
    .B(_01778_),
    .Y(_01783_)
  );
  INVX1 _08452_ (
    .A(_01783_),
    .Y(_01784_)
  );
  NAND2X1 _08453_ (
    .A(_01747_),
    .B(_01763_),
    .Y(_01785_)
  );
  AOI21X1 _08454_ (
    .A(_01747_),
    .B(_01763_),
    .C(_01784_),
    .Y(_01786_)
  );
  OAI21X1 _08455_ (
    .A(_01746_),
    .B(_01762_),
    .C(_01783_),
    .Y(_01787_)
  );
  XNOR2X1 _08456_ (
    .A(_01784_),
    .B(_01785_),
    .Y(_01788_)
  );
  XNOR2X1 _08457_ (
    .A(_01783_),
    .B(_01785_),
    .Y(_01789_)
  );
  XOR2X1 _08458_ (
    .A( execution_unit_0.alu_0.alu_shift_14_ ),
    .B(_01386_),
    .Y(_01790_)
  );
  NOR2X1 _08459_ (
    .A(_01622_),
    .B(_01790_),
    .Y(_01791_)
  );
  OAI21X1 _08460_ (
    .A(_01899_),
    .B(_01371_),
    .C( execution_unit_0.alu_0.op_dst_15_ ),
    .Y(_01792_)
  );
  NOR2X1 _08461_ (
    .A(_01790_),
    .B(_01792_),
    .Y(_01793_)
  );
  NAND2X1 _08462_ (
    .A( execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01791_),
    .Y(_01794_)
  );
  OAI21X1 _08463_ (
    .A(_01622_),
    .B(_01790_),
    .C(_01792_),
    .Y(_01795_)
  );
  XOR2X1 _08464_ (
    .A( execution_unit_0.alu_0.alu_shift_13_ ),
    .B(_01386_),
    .Y(_01796_)
  );
  NOR2X1 _08465_ (
    .A(_01622_),
    .B(_01796_),
    .Y(_01797_)
  );
  AND2X1 _08466_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01623_),
    .Y(_01798_)
  );
  AND2X1 _08467_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01797_),
    .Y(_01799_)
  );
  NAND2X1 _08468_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01797_),
    .Y(_01800_)
  );
  NOR2X1 _08469_ (
    .A(_01797_),
    .B(_01798_),
    .Y(_01801_)
  );
  NOR2X1 _08470_ (
    .A(_01799_),
    .B(_01801_),
    .Y(_01802_)
  );
  OAI21X1 _08471_ (
    .A(_01797_),
    .B(_01798_),
    .C(_01800_),
    .Y(_01803_)
  );
  AOI21X1 _08472_ (
    .A(_01777_),
    .B(_01787_),
    .C(_01803_),
    .Y(_01804_)
  );
  OAI21X1 _08473_ (
    .A(_01776_),
    .B(_01786_),
    .C(_01802_),
    .Y(_01805_)
  );
  OAI21X1 _08474_ (
    .A(_01799_),
    .B(_01804_),
    .C(_01795_),
    .Y(_01806_)
  );
  AND2X1 _08475_ (
    .A(_01794_),
    .B(_01806_),
    .Y(_01807_)
  );
  OAI21X1 _08476_ (
    .A(_01790_),
    .B(_01792_),
    .C(_01806_),
    .Y(_01808_)
  );
  NOR3X1 _08477_ (
    .A(_01776_),
    .B(_01786_),
    .C(_01802_),
    .Y(_01809_)
  );
  NAND3X1 _08478_ (
    .A(_01777_),
    .B(_01787_),
    .C(_01803_),
    .Y(_01810_)
  );
  NOR2X1 _08479_ (
    .A(_01804_),
    .B(_01809_),
    .Y(_01811_)
  );
  AOI21X1 _08480_ (
    .A(_01805_),
    .B(_01810_),
    .C(_01788_),
    .Y(_01812_)
  );
  OAI21X1 _08481_ (
    .A(_01804_),
    .B(_01809_),
    .C(_01789_),
    .Y(_01813_)
  );
  AND2X1 _08482_ (
    .A(_01794_),
    .B(_01795_),
    .Y(_01814_)
  );
  OAI21X1 _08483_ (
    .A(_01790_),
    .B(_01792_),
    .C(_01795_),
    .Y(_01815_)
  );
  NOR3X1 _08484_ (
    .A(_01799_),
    .B(_01804_),
    .C(_01814_),
    .Y(_01816_)
  );
  NAND3X1 _08485_ (
    .A(_01800_),
    .B(_01805_),
    .C(_01815_),
    .Y(_01817_)
  );
  AOI21X1 _08486_ (
    .A(_01800_),
    .B(_01805_),
    .C(_01815_),
    .Y(_01818_)
  );
  OAI21X1 _08487_ (
    .A(_01799_),
    .B(_01804_),
    .C(_01814_),
    .Y(_01819_)
  );
  NOR3X1 _08488_ (
    .A(_01812_),
    .B(_01816_),
    .C(_01818_),
    .Y(_01820_)
  );
  NAND3X1 _08489_ (
    .A(_01813_),
    .B(_01817_),
    .C(_01819_),
    .Y(_01821_)
  );
  AOI21X1 _08490_ (
    .A(_01807_),
    .B(_01821_),
    .C(_01788_),
    .Y(_01822_)
  );
  OAI21X1 _08491_ (
    .A(_01808_),
    .B(_01820_),
    .C(_01789_),
    .Y(_01823_)
  );
  NOR3X1 _08492_ (
    .A(_01789_),
    .B(_01808_),
    .C(_01820_),
    .Y(_01824_)
  );
  NOR3X1 _08493_ (
    .A(_01368_),
    .B(_01822_),
    .C(_01824_),
    .Y(_01825_)
  );
  NOR2X1 _08494_ (
    .A(_01365_),
    .B(_01784_),
    .Y(_01826_)
  );
  NAND2X1 _08495_ (
    .A(_01400_),
    .B(_01775_),
    .Y(_01827_)
  );
  AOI22X1 _08496_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_13_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01828_)
  );
  NAND3X1 _08497_ (
    .A(_01612_),
    .B(_01827_),
    .C(_01828_),
    .Y(_01829_)
  );
  AOI21X1 _08498_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01776_),
    .C(_01829_),
    .Y(_01830_)
  );
  OAI21X1 _08499_ (
    .A(_01364_),
    .B(_01778_),
    .C(_01830_),
    .Y(_01831_)
  );
  OAI21X1 _08500_ (
    .A(_01826_),
    .B(_01831_),
    .C(_01373_),
    .Y(_01832_)
  );
  OAI22X1 _08501_ (
    .A(_01373_),
    .B(_01782_),
    .C(_01825_),
    .D(_01832_),
    .Y( execution_unit_0.alu_0.alu_out_13_ )
  );
  OAI22X1 _08502_ (
    .A(_01385_),
    .B(_01777_),
    .C(_01778_),
    .D(_01748_),
    .Y(_01833_)
  );
  INVX1 _08503_ (
    .A(_01833_),
    .Y(_01834_)
  );
  OAI21X1 _08504_ (
    .A(_01752_),
    .B(_01779_),
    .C(_01834_),
    .Y(_01835_)
  );
  AOI21X1 _08505_ (
    .A(_01384_),
    .B(_01797_),
    .C(_01798_),
    .Y(_01836_)
  );
  AOI21X1 _08506_ (
    .A(_01384_),
    .B(_01799_),
    .C(_01836_),
    .Y(_01837_)
  );
  NAND2X1 _08507_ (
    .A(_01835_),
    .B(_01837_),
    .Y(_01838_)
  );
  XOR2X1 _08508_ (
    .A(_01835_),
    .B(_01837_),
    .Y( dbg_0.UNUSED_eu_mab_14_ )
  );
  OAI21X1 _08509_ (
    .A(_01807_),
    .B(_01813_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01839_)
  );
  AOI21X1 _08510_ (
    .A(_01811_),
    .B(_01823_),
    .C(_01839_),
    .Y(_01840_)
  );
  OAI21X1 _08511_ (
    .A(_01797_),
    .B(_01798_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01841_)
  );
  AOI22X1 _08512_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C( execution_unit_0.alu_0.alu_shift_14_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01842_)
  );
  AOI22X1 _08513_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C(_01400_),
    .D(_01797_),
    .Y(_01843_)
  );
  OAI21X1 _08514_ (
    .A(_01363_),
    .B(_01800_),
    .C(_01843_),
    .Y(_01844_)
  );
  AOI21X1 _08515_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01802_),
    .C(_01844_),
    .Y(_01845_)
  );
  NAND3X1 _08516_ (
    .A(_01841_),
    .B(_01842_),
    .C(_01845_),
    .Y(_01846_)
  );
  OAI21X1 _08517_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01846_),
    .C(_01373_),
    .Y(_01847_)
  );
  AND2X1 _08518_ (
    .A(_01781_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_01848_)
  );
  NAND2X1 _08519_ (
    .A(_01781_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_01849_)
  );
  OAI21X1 _08520_ (
    .A(_01781_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .C(_01374_),
    .Y(_01850_)
  );
  OAI22X1 _08521_ (
    .A(_01840_),
    .B(_01847_),
    .C(_01848_),
    .D(_01850_),
    .Y( execution_unit_0.alu_0.alu_out_14_ )
  );
  NAND2X1 _08522_ (
    .A(_01384_),
    .B(_01791_),
    .Y(_01851_)
  );
  AOI22X1 _08523_ (
    .A(_01384_),
    .B(_01793_),
    .C(_01851_),
    .D(_01792_),
    .Y(_01852_)
  );
  OAI21X1 _08524_ (
    .A(_01385_),
    .B(_01800_),
    .C(_01838_),
    .Y(_01853_)
  );
  XOR2X1 _08525_ (
    .A(_01852_),
    .B(_01853_),
    .Y( dbg_0.UNUSED_eu_mab_15_ )
  );
  INVX1 _08526_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_01854_)
  );
  XNOR2X1 _08527_ (
    .A(_01849_),
    .B( dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_01855_)
  );
  NOR2X1 _08528_ (
    .A(_01373_),
    .B(_01855_),
    .Y(_01856_)
  );
  AND2X1 _08529_ (
    .A(_01400_),
    .B(_01791_),
    .Y(_01857_)
  );
  OAI21X1 _08530_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01858_)
  );
  OAI21X1 _08531_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01857_),
    .C(_01795_),
    .Y(_01859_)
  );
  OAI22X1 _08532_ (
    .A(_01366_),
    .B(_01609_),
    .C(_01794_),
    .D(_01363_),
    .Y(_01860_)
  );
  AOI21X1 _08533_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01814_),
    .C(_01860_),
    .Y(_01861_)
  );
  NAND3X1 _08534_ (
    .A(_01858_),
    .B(_01859_),
    .C(_01861_),
    .Y(_01862_)
  );
  INVX1 _08535_ (
    .A(_01862_),
    .Y(_01863_)
  );
  OAI21X1 _08536_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01863_),
    .C(_01373_),
    .Y(_01864_)
  );
  OAI22X1 _08537_ (
    .A(_01807_),
    .B(_01812_),
    .C(_01816_),
    .D(_01818_),
    .Y(_01865_)
  );
  NOR2X1 _08538_ (
    .A(_01368_),
    .B(_01820_),
    .Y(_01866_)
  );
  AOI21X1 _08539_ (
    .A(_01865_),
    .B(_01866_),
    .C(_01864_),
    .Y(_01867_)
  );
  NOR2X1 _08540_ (
    .A(_01856_),
    .B(_01867_),
    .Y( execution_unit_0.alu_0.alu_out_15_ )
  );
  NAND2X1 _08541_ (
    .A(_01371_),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_01868_)
  );
  OAI21X1 _08542_ (
    .A(_01371_),
    .B(_01619_),
    .C(_01868_),
    .Y( execution_unit_0.alu_0.N )
  );
  NAND3X1 _08543_ (
    .A(_01651_),
    .B(_01704_),
    .C(_01742_),
    .Y(_01869_)
  );
  OR2X1 _08544_ (
    .A( execution_unit_0.alu_0.alu_out_10_ ),
    .B(_01869_),
    .Y(_01870_)
  );
  NOR2X1 _08545_ (
    .A( execution_unit_0.alu_0.alu_out_12_ ),
    .B(_01870_),
    .Y(_01871_)
  );
  OAI21X1 _08546_ (
    .A(_01856_),
    .B(_01867_),
    .C(_01871_),
    .Y(_01872_)
  );
  NOR3X1 _08547_ (
    .A( execution_unit_0.alu_0.alu_out_13_ ),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .C(_01872_),
    .Y(_01873_)
  );
  OR2X1 _08548_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_01874_)
  );
  NOR2X1 _08549_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_01874_),
    .Y(_01875_)
  );
  NOR2X1 _08550_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_01876_)
  );
  NAND3X1 _08551_ (
    .A(_01619_),
    .B(_01875_),
    .C(_01876_),
    .Y(_01877_)
  );
  NOR3X1 _08552_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .C(_01877_),
    .Y(_01878_)
  );
  OAI21X1 _08553_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01873_),
    .C(_01878_),
    .Y(_01879_)
  );
  INVX1 _08554_ (
    .A(_01879_),
    .Y( execution_unit_0.alu_0.Z )
  );
  NAND2X1 _08555_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01387_),
    .Y(_01880_)
  );
  NOR2X1 _08556_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B( execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01881_)
  );
  NOR2X1 _08557_ (
    .A(_01879_),
    .B(_01881_),
    .Y(_01882_)
  );
  AOI22X1 _08558_ (
    .A(_01384_),
    .B(_01793_),
    .C(_01852_),
    .D(_01853_),
    .Y(_01883_)
  );
  OAI21X1 _08559_ (
    .A(_01849_),
    .B(_01854_),
    .C(_01883_),
    .Y(_01884_)
  );
  OAI21X1 _08560_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01372_),
    .C(_01884_),
    .Y(_01885_)
  );
  AOI21X1 _08561_ (
    .A(_01807_),
    .B(_01821_),
    .C(_01469_),
    .Y(_01886_)
  );
  OAI21X1 _08562_ (
    .A(_01807_),
    .B(_01821_),
    .C(_01886_),
    .Y(_01887_)
  );
  AOI21X1 _08563_ (
    .A(_01885_),
    .B(_01887_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_01888_)
  );
  OAI21X1 _08564_ (
    .A(_01371_),
    .B(_01651_),
    .C(_01881_),
    .Y(_01889_)
  );
  OAI21X1 _08565_ (
    .A(_01888_),
    .B(_01889_),
    .C(_01366_),
    .Y(_01890_)
  );
  OAI21X1 _08566_ (
    .A(_01882_),
    .B(_01890_),
    .C(_01880_),
    .Y( execution_unit_0.alu_0.alu_stat_0_ )
  );
  NOR2X1 _08567_ (
    .A(_01554_),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01891_)
  );
  OAI21X1 _08568_ (
    .A(_01555_),
    .B(_01619_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_01892_)
  );
  MUX2X1 _08569_ (
    .A(_01795_),
    .B(_01794_),
    .S( execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_01893_)
  );
  OAI22X1 _08570_ (
    .A(_01891_),
    .B(_01892_),
    .C(_01893_),
    .D( execution_unit_0.alu_0.inst_bw ),
    .Y(_01894_)
  );
  NOR2X1 _08571_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01794_),
    .Y(_01895_)
  );
  OAI21X1 _08572_ (
    .A(_01371_),
    .B(_01554_),
    .C( execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01896_)
  );
  NOR2X1 _08573_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01897_)
  );
  OAI21X1 _08574_ (
    .A(_01895_),
    .B(_01896_),
    .C(_01897_),
    .Y(_01898_)
  );
  AOI21X1 _08575_ (
    .A(_01365_),
    .B(_01894_),
    .C(_01898_),
    .Y( execution_unit_0.alu_0.alu_stat_3_ )
  );
  AND2X1 _08576_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .B( execution_unit_0.alu_0.inst_alu_9_ ),
    .Y( execution_unit_0.alu_0.alu_stat_wr_0_ )
  );
  INVX1 _08577_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_03094_)
  );
  INVX1 _08578_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_03095_)
  );
  INVX1 _08579_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_03096_)
  );
  INVX1 _08580_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_03097_)
  );
  INVX1 _08581_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_03098_)
  );
  INVX1 _08582_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_03099_)
  );
  INVX1 _08583_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_03100_)
  );
  INVX1 _08584_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_03101_)
  );
  INVX1 _08585_ (
    .A( execution_unit_0.register_file_0.r4_10_ ),
    .Y(_03102_)
  );
  INVX1 _08586_ (
    .A( execution_unit_0.register_file_0.r4_1_ ),
    .Y(_03103_)
  );
  INVX1 _08587_ (
    .A( execution_unit_0.reg_sp_wr ),
    .Y(_03104_)
  );
  INVX1 _08588_ (
    .A( execution_unit_0.reg_sr_clr ),
    .Y(_03105_)
  );
  INVX1 _08589_ (
    .A( execution_unit_0.inst_src_1_ ),
    .Y(_03106_)
  );
  INVX1 _08590_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_03107_)
  );
  INVX1 _08591_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .Y(_03108_)
  );
  INVX1 _08592_ (
    .A( execution_unit_0.register_file_0.r2_4_ ),
    .Y(_03109_)
  );
  INVX1 _08593_ (
    .A( execution_unit_0.alu_0.alu_stat_3_ ),
    .Y(_03110_)
  );
  INVX1 _08594_ (
    .A(_06327_),
    .Y(_01901_)
  );
  AND2X1 _08595_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_13_ ),
    .Y(_03111_)
  );
  AND2X1 _08596_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_11_ ),
    .Y(_03112_)
  );
  NOR2X1 _08597_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_03106_),
    .Y(_03113_)
  );
  AND2X1 _08598_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_9_ ),
    .Y(_03114_)
  );
  AND2X1 _08599_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_10_ ),
    .Y(_03115_)
  );
  AND2X1 _08600_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_8_ ),
    .Y(_03116_)
  );
  AND2X1 _08601_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_0_ ),
    .Y(_03117_)
  );
  NAND2X1 _08602_ (
    .A( dbg_0.UNUSED_pc_14_ ),
    .B(_03117_),
    .Y(_03118_)
  );
  AND2X1 _08603_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_15_ ),
    .Y(_03119_)
  );
  AND2X1 _08604_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_7_ ),
    .Y(_03120_)
  );
  NAND2X1 _08605_ (
    .A( execution_unit_0.register_file_0.r7_14_ ),
    .B(_03120_),
    .Y(_03121_)
  );
  AND2X1 _08606_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_5_ ),
    .Y(_03122_)
  );
  AND2X1 _08607_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_14_ ),
    .Y(_03123_)
  );
  AND2X1 _08608_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_6_ ),
    .Y(_03124_)
  );
  AND2X1 _08609_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_12_ ),
    .Y(_03125_)
  );
  AND2X1 _08610_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_4_ ),
    .Y(_03126_)
  );
  NAND2X1 _08611_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_4_ ),
    .Y(_03127_)
  );
  AND2X1 _08612_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_3_ ),
    .Y(_03128_)
  );
  AOI22X1 _08613_ (
    .A( execution_unit_0.register_file_0.r13_14_ ),
    .B(_03111_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_14_ ),
    .Y(_03129_)
  );
  AOI22X1 _08614_ (
    .A( execution_unit_0.register_file_0.r5_14_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_14_ ),
    .Y(_03130_)
  );
  AOI22X1 _08615_ (
    .A( execution_unit_0.register_file_0.r1_14_ ),
    .B(_03113_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_14_ ),
    .Y(_03131_)
  );
  NAND2X1 _08616_ (
    .A(_03130_),
    .B(_03131_),
    .Y(_03132_)
  );
  AOI21X1 _08617_ (
    .A( execution_unit_0.register_file_0.r6_14_ ),
    .B(_03124_),
    .C(_03132_),
    .Y(_03133_)
  );
  NAND3X1 _08618_ (
    .A(_03118_),
    .B(_03121_),
    .C(_03129_),
    .Y(_03134_)
  );
  AOI22X1 _08619_ (
    .A( execution_unit_0.register_file_0.r11_14_ ),
    .B(_03112_),
    .C(_03114_),
    .D( execution_unit_0.register_file_0.r9_14_ ),
    .Y(_03135_)
  );
  AOI22X1 _08620_ (
    .A( execution_unit_0.register_file_0.r10_14_ ),
    .B(_03115_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_03136_)
  );
  AOI22X1 _08621_ (
    .A( execution_unit_0.register_file_0.r8_14_ ),
    .B(_03116_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_14_ ),
    .Y(_03137_)
  );
  NAND3X1 _08622_ (
    .A(_03135_),
    .B(_03136_),
    .C(_03137_),
    .Y(_03138_)
  );
  NOR2X1 _08623_ (
    .A(_03134_),
    .B(_03138_),
    .Y(_03139_)
  );
  NAND2X1 _08624_ (
    .A(_03133_),
    .B(_03139_),
    .Y( execution_unit_0.reg_src_14_ )
  );
  INVX1 _08625_ (
    .A( execution_unit_0.reg_src_14_ ),
    .Y(_03140_)
  );
  AOI22X1 _08626_ (
    .A( execution_unit_0.register_file_0.r5_13_ ),
    .B(_03122_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_13_ ),
    .Y(_03141_)
  );
  NAND2X1 _08627_ (
    .A( execution_unit_0.register_file_0.r14_13_ ),
    .B(_03123_),
    .Y(_03142_)
  );
  AOI22X1 _08628_ (
    .A( execution_unit_0.register_file_0.r13_13_ ),
    .B(_03111_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_13_ ),
    .Y(_03143_)
  );
  AOI22X1 _08629_ (
    .A( execution_unit_0.register_file_0.r8_13_ ),
    .B(_03116_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_13_ ),
    .Y(_03144_)
  );
  AOI22X1 _08630_ (
    .A( execution_unit_0.register_file_0.r9_13_ ),
    .B(_03114_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_13_ ),
    .Y(_03145_)
  );
  NAND2X1 _08631_ (
    .A(_03142_),
    .B(_03145_),
    .Y(_03146_)
  );
  AOI21X1 _08632_ (
    .A( execution_unit_0.register_file_0.r7_13_ ),
    .B(_03120_),
    .C(_03146_),
    .Y(_03147_)
  );
  AND2X1 _08633_ (
    .A(_03143_),
    .B(_03144_),
    .Y(_03148_)
  );
  AOI22X1 _08634_ (
    .A( execution_unit_0.register_file_0.r11_13_ ),
    .B(_03112_),
    .C(_03115_),
    .D( execution_unit_0.register_file_0.r10_13_ ),
    .Y(_03149_)
  );
  AOI22X1 _08635_ (
    .A( dbg_0.UNUSED_pc_13_ ),
    .B(_03117_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_13_ ),
    .Y(_03150_)
  );
  NAND3X1 _08636_ (
    .A(_03141_),
    .B(_03149_),
    .C(_03150_),
    .Y(_03151_)
  );
  AOI21X1 _08637_ (
    .A( execution_unit_0.register_file_0.r1_13_ ),
    .B(_03113_),
    .C(_03151_),
    .Y(_03152_)
  );
  NAND3X1 _08638_ (
    .A(_03147_),
    .B(_03148_),
    .C(_03152_),
    .Y( execution_unit_0.reg_src_13_ )
  );
  INVX1 _08639_ (
    .A( execution_unit_0.reg_src_13_ ),
    .Y(_03153_)
  );
  AOI22X1 _08640_ (
    .A( execution_unit_0.register_file_0.r13_12_ ),
    .B(_03111_),
    .C(_03115_),
    .D( execution_unit_0.register_file_0.r10_12_ ),
    .Y(_03154_)
  );
  AOI22X1 _08641_ (
    .A( execution_unit_0.register_file_0.r9_12_ ),
    .B(_03114_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_12_ ),
    .Y(_03155_)
  );
  NAND2X1 _08642_ (
    .A(_03154_),
    .B(_03155_),
    .Y(_03156_)
  );
  AOI22X1 _08643_ (
    .A( execution_unit_0.register_file_0.r11_12_ ),
    .B(_03112_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_12_ ),
    .Y(_03157_)
  );
  AOI22X1 _08644_ (
    .A( execution_unit_0.register_file_0.r8_12_ ),
    .B(_03116_),
    .C(_03117_),
    .D( dbg_0.UNUSED_pc_12_ ),
    .Y(_03158_)
  );
  NAND2X1 _08645_ (
    .A(_03157_),
    .B(_03158_),
    .Y(_03159_)
  );
  NOR2X1 _08646_ (
    .A(_03156_),
    .B(_03159_),
    .Y(_03160_)
  );
  NAND2X1 _08647_ (
    .A( execution_unit_0.register_file_0.r7_12_ ),
    .B(_03120_),
    .Y(_03161_)
  );
  AOI22X1 _08648_ (
    .A( execution_unit_0.register_file_0.r1_12_ ),
    .B(_03113_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_12_ ),
    .Y(_03162_)
  );
  NAND2X1 _08649_ (
    .A(_03161_),
    .B(_03162_),
    .Y(_03163_)
  );
  AOI22X1 _08650_ (
    .A( execution_unit_0.register_file_0.r5_12_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_12_ ),
    .Y(_03164_)
  );
  AOI22X1 _08651_ (
    .A( execution_unit_0.register_file_0.r15_12_ ),
    .B(_03119_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_12_ ),
    .Y(_03165_)
  );
  NAND2X1 _08652_ (
    .A(_03164_),
    .B(_03165_),
    .Y(_03166_)
  );
  NOR2X1 _08653_ (
    .A(_03163_),
    .B(_03166_),
    .Y(_03167_)
  );
  NAND2X1 _08654_ (
    .A(_03160_),
    .B(_03167_),
    .Y( execution_unit_0.reg_src_12_ )
  );
  INVX1 _08655_ (
    .A( execution_unit_0.reg_src_12_ ),
    .Y(_03168_)
  );
  NAND2X1 _08656_ (
    .A( dbg_0.UNUSED_pc_11_ ),
    .B(_03117_),
    .Y(_03169_)
  );
  NAND2X1 _08657_ (
    .A( execution_unit_0.register_file_0.r7_11_ ),
    .B(_03120_),
    .Y(_03170_)
  );
  AOI22X1 _08658_ (
    .A( execution_unit_0.register_file_0.r10_11_ ),
    .B(_03115_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_11_ ),
    .Y(_03171_)
  );
  AOI22X1 _08659_ (
    .A( execution_unit_0.register_file_0.r11_11_ ),
    .B(_03112_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_11_ ),
    .Y(_03172_)
  );
  AOI22X1 _08660_ (
    .A( execution_unit_0.register_file_0.r13_11_ ),
    .B(_03111_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_11_ ),
    .Y(_03173_)
  );
  AOI22X1 _08661_ (
    .A( execution_unit_0.register_file_0.r5_11_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_11_ ),
    .Y(_03174_)
  );
  AOI22X1 _08662_ (
    .A( execution_unit_0.register_file_0.r6_11_ ),
    .B(_03124_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_11_ ),
    .Y(_03175_)
  );
  NAND2X1 _08663_ (
    .A(_03174_),
    .B(_03175_),
    .Y(_03176_)
  );
  AOI21X1 _08664_ (
    .A( execution_unit_0.register_file_0.r1_11_ ),
    .B(_03113_),
    .C(_03176_),
    .Y(_03177_)
  );
  NAND3X1 _08665_ (
    .A(_03169_),
    .B(_03170_),
    .C(_03173_),
    .Y(_03178_)
  );
  AOI22X1 _08666_ (
    .A( execution_unit_0.register_file_0.r9_11_ ),
    .B(_03114_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_11_ ),
    .Y(_03179_)
  );
  NAND3X1 _08667_ (
    .A(_03171_),
    .B(_03172_),
    .C(_03179_),
    .Y(_03180_)
  );
  NOR2X1 _08668_ (
    .A(_03178_),
    .B(_03180_),
    .Y(_03181_)
  );
  NAND2X1 _08669_ (
    .A(_03177_),
    .B(_03181_),
    .Y( execution_unit_0.reg_src_11_ )
  );
  INVX1 _08670_ (
    .A( execution_unit_0.reg_src_11_ ),
    .Y(_03182_)
  );
  NAND2X1 _08671_ (
    .A( execution_unit_0.register_file_0.r11_10_ ),
    .B(_03112_),
    .Y(_03183_)
  );
  AOI22X1 _08672_ (
    .A( execution_unit_0.register_file_0.r8_10_ ),
    .B(_03116_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_10_ ),
    .Y(_03184_)
  );
  OAI21X1 _08673_ (
    .A(_03102_),
    .B(_03127_),
    .C(_03184_),
    .Y(_03185_)
  );
  AOI22X1 _08674_ (
    .A( execution_unit_0.register_file_0.r1_10_ ),
    .B(_03113_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_10_ ),
    .Y(_03186_)
  );
  AOI22X1 _08675_ (
    .A( execution_unit_0.register_file_0.r10_10_ ),
    .B(_03115_),
    .C(_03122_),
    .D( execution_unit_0.register_file_0.r5_10_ ),
    .Y(_03187_)
  );
  AOI22X1 _08676_ (
    .A( execution_unit_0.register_file_0.r9_10_ ),
    .B(_03114_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_10_ ),
    .Y(_03188_)
  );
  NAND3X1 _08677_ (
    .A(_03186_),
    .B(_03187_),
    .C(_03188_),
    .Y(_03189_)
  );
  AOI21X1 _08678_ (
    .A( execution_unit_0.register_file_0.r13_10_ ),
    .B(_03111_),
    .C(_03189_),
    .Y(_03190_)
  );
  AOI22X1 _08679_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .B(_03117_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_10_ ),
    .Y(_03191_)
  );
  AOI22X1 _08680_ (
    .A( execution_unit_0.register_file_0.r15_10_ ),
    .B(_03119_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_10_ ),
    .Y(_03192_)
  );
  NAND2X1 _08681_ (
    .A(_03183_),
    .B(_03192_),
    .Y(_03193_)
  );
  NOR2X1 _08682_ (
    .A(_03185_),
    .B(_03193_),
    .Y(_03194_)
  );
  NAND3X1 _08683_ (
    .A(_03190_),
    .B(_03191_),
    .C(_03194_),
    .Y( execution_unit_0.reg_src_10_ )
  );
  INVX1 _08684_ (
    .A( execution_unit_0.reg_src_10_ ),
    .Y(_03195_)
  );
  NAND2X1 _08685_ (
    .A( execution_unit_0.register_file_0.r1_9_ ),
    .B(_03113_),
    .Y(_03196_)
  );
  NAND2X1 _08686_ (
    .A( dbg_0.UNUSED_pc_9_ ),
    .B(_03117_),
    .Y(_03197_)
  );
  AOI22X1 _08687_ (
    .A( execution_unit_0.register_file_0.r9_9_ ),
    .B(_03114_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_9_ ),
    .Y(_03198_)
  );
  AOI22X1 _08688_ (
    .A( execution_unit_0.register_file_0.r10_9_ ),
    .B(_03115_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_9_ ),
    .Y(_03199_)
  );
  AOI22X1 _08689_ (
    .A( execution_unit_0.register_file_0.r11_9_ ),
    .B(_03112_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_9_ ),
    .Y(_03200_)
  );
  NAND3X1 _08690_ (
    .A(_03198_),
    .B(_03199_),
    .C(_03200_),
    .Y(_03201_)
  );
  AOI21X1 _08691_ (
    .A( execution_unit_0.register_file_0.r7_9_ ),
    .B(_03120_),
    .C(_03201_),
    .Y(_03202_)
  );
  AOI22X1 _08692_ (
    .A( execution_unit_0.register_file_0.r13_9_ ),
    .B(_03111_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_9_ ),
    .Y(_03203_)
  );
  AOI22X1 _08693_ (
    .A( execution_unit_0.register_file_0.r5_9_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_9_ ),
    .Y(_03204_)
  );
  NAND2X1 _08694_ (
    .A(_03196_),
    .B(_03204_),
    .Y(_03205_)
  );
  AOI22X1 _08695_ (
    .A( execution_unit_0.register_file_0.r6_9_ ),
    .B(_03124_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_9_ ),
    .Y(_03206_)
  );
  NAND2X1 _08696_ (
    .A(_03197_),
    .B(_03206_),
    .Y(_03207_)
  );
  NOR2X1 _08697_ (
    .A(_03205_),
    .B(_03207_),
    .Y(_03208_)
  );
  NAND3X1 _08698_ (
    .A(_03202_),
    .B(_03203_),
    .C(_03208_),
    .Y( execution_unit_0.reg_src_9_ )
  );
  INVX1 _08699_ (
    .A( execution_unit_0.reg_src_9_ ),
    .Y(_03209_)
  );
  AOI22X1 _08700_ (
    .A( execution_unit_0.register_file_0.r10_8_ ),
    .B(_03115_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_8_ ),
    .Y(_03210_)
  );
  AOI22X1 _08701_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .B(_03117_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_8_ ),
    .Y(_03211_)
  );
  AOI22X1 _08702_ (
    .A( execution_unit_0.register_file_0.r11_8_ ),
    .B(_03112_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_8_ ),
    .Y(_03212_)
  );
  AOI22X1 _08703_ (
    .A( execution_unit_0.register_file_0.r13_8_ ),
    .B(_03111_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_8_ ),
    .Y(_03213_)
  );
  AND2X1 _08704_ (
    .A(_03212_),
    .B(_03213_),
    .Y(_03214_)
  );
  NAND3X1 _08705_ (
    .A(_03210_),
    .B(_03211_),
    .C(_03214_),
    .Y(_03215_)
  );
  OR2X1 _08706_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .Y(_03216_)
  );
  AOI22X1 _08707_ (
    .A( execution_unit_0.register_file_0.r7_8_ ),
    .B(_03120_),
    .C(_03216_),
    .D( execution_unit_0.alu_0.status_3_ ),
    .Y(_03217_)
  );
  AOI22X1 _08708_ (
    .A( execution_unit_0.register_file_0.r5_8_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_8_ ),
    .Y(_03218_)
  );
  AOI22X1 _08709_ (
    .A( execution_unit_0.register_file_0.r14_8_ ),
    .B(_03123_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_8_ ),
    .Y(_03219_)
  );
  AOI22X1 _08710_ (
    .A( execution_unit_0.register_file_0.r1_8_ ),
    .B(_03113_),
    .C(_03114_),
    .D( execution_unit_0.register_file_0.r9_8_ ),
    .Y(_03220_)
  );
  AND2X1 _08711_ (
    .A(_03219_),
    .B(_03220_),
    .Y(_03221_)
  );
  NAND3X1 _08712_ (
    .A(_03217_),
    .B(_03218_),
    .C(_03221_),
    .Y(_03222_)
  );
  NOR2X1 _08713_ (
    .A(_03215_),
    .B(_03222_),
    .Y(_03223_)
  );
  INVX1 _08714_ (
    .A(_03223_),
    .Y( execution_unit_0.reg_src_8_ )
  );
  AOI22X1 _08715_ (
    .A( execution_unit_0.register_file_0.r4_7_ ),
    .B(_03126_),
    .C(_03216_),
    .D( clock_module_0.scg1 ),
    .Y(_03224_)
  );
  AOI22X1 _08716_ (
    .A( execution_unit_0.register_file_0.r10_7_ ),
    .B(_03115_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_7_ ),
    .Y(_03225_)
  );
  AOI22X1 _08717_ (
    .A( execution_unit_0.register_file_0.r6_7_ ),
    .B(_03124_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_7_ ),
    .Y(_03226_)
  );
  AOI22X1 _08718_ (
    .A( execution_unit_0.register_file_0.r8_7_ ),
    .B(_03116_),
    .C(_03122_),
    .D( execution_unit_0.register_file_0.r5_7_ ),
    .Y(_03227_)
  );
  AND2X1 _08719_ (
    .A(_03226_),
    .B(_03227_),
    .Y(_03228_)
  );
  NAND3X1 _08720_ (
    .A(_03224_),
    .B(_03225_),
    .C(_03228_),
    .Y(_03229_)
  );
  AOI22X1 _08721_ (
    .A( execution_unit_0.register_file_0.r11_7_ ),
    .B(_03112_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_7_ ),
    .Y(_03230_)
  );
  AOI22X1 _08722_ (
    .A( execution_unit_0.register_file_0.r13_7_ ),
    .B(_03111_),
    .C(_03114_),
    .D( execution_unit_0.register_file_0.r9_7_ ),
    .Y(_03231_)
  );
  AOI22X1 _08723_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .B(_03117_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_7_ ),
    .Y(_03232_)
  );
  AOI22X1 _08724_ (
    .A( execution_unit_0.register_file_0.r1_7_ ),
    .B(_03113_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_7_ ),
    .Y(_03233_)
  );
  AND2X1 _08725_ (
    .A(_03232_),
    .B(_03233_),
    .Y(_03234_)
  );
  NAND3X1 _08726_ (
    .A(_03230_),
    .B(_03231_),
    .C(_03234_),
    .Y(_03235_)
  );
  NOR2X1 _08727_ (
    .A(_03229_),
    .B(_03235_),
    .Y(_03236_)
  );
  INVX1 _08728_ (
    .A(_03236_),
    .Y( execution_unit_0.reg_src_7_ )
  );
  AOI22X1 _08729_ (
    .A( execution_unit_0.register_file_0.r9_6_ ),
    .B(_03114_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_6_ ),
    .Y(_03237_)
  );
  AOI22X1 _08730_ (
    .A( execution_unit_0.register_file_0.r1_6_ ),
    .B(_03113_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_6_ ),
    .Y(_03238_)
  );
  AOI22X1 _08731_ (
    .A( execution_unit_0.register_file_0.r13_6_ ),
    .B(_03111_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_6_ ),
    .Y(_03239_)
  );
  AOI22X1 _08732_ (
    .A( execution_unit_0.register_file_0.r10_6_ ),
    .B(_03115_),
    .C(_03122_),
    .D( execution_unit_0.register_file_0.r5_6_ ),
    .Y(_03240_)
  );
  AND2X1 _08733_ (
    .A(_03239_),
    .B(_03240_),
    .Y(_03241_)
  );
  NAND3X1 _08734_ (
    .A(_03237_),
    .B(_03238_),
    .C(_03241_),
    .Y(_03242_)
  );
  AOI22X1 _08735_ (
    .A( execution_unit_0.register_file_0.r15_6_ ),
    .B(_03119_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_6_ ),
    .Y(_03243_)
  );
  INVX1 _08736_ (
    .A(_03243_),
    .Y(_03244_)
  );
  AOI21X1 _08737_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B(_03117_),
    .C(_03244_),
    .Y(_03245_)
  );
  AOI22X1 _08738_ (
    .A( execution_unit_0.register_file_0.r14_6_ ),
    .B(_03123_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_6_ ),
    .Y(_03246_)
  );
  AOI22X1 _08739_ (
    .A( execution_unit_0.register_file_0.r11_6_ ),
    .B(_03112_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_6_ ),
    .Y(_03247_)
  );
  NAND3X1 _08740_ (
    .A(_03245_),
    .B(_03246_),
    .C(_03247_),
    .Y(_03248_)
  );
  OR2X1 _08741_ (
    .A(_03242_),
    .B(_03248_),
    .Y( execution_unit_0.reg_src_6_ )
  );
  INVX1 _08742_ (
    .A( execution_unit_0.reg_src_6_ ),
    .Y(_03249_)
  );
  AOI22X1 _08743_ (
    .A( execution_unit_0.register_file_0.r13_5_ ),
    .B(_03111_),
    .C(_03122_),
    .D( execution_unit_0.register_file_0.r5_5_ ),
    .Y(_03250_)
  );
  AOI22X1 _08744_ (
    .A( execution_unit_0.register_file_0.r15_5_ ),
    .B(_03119_),
    .C(_03216_),
    .D( clock_module_0.oscoff ),
    .Y(_03251_)
  );
  NAND2X1 _08745_ (
    .A(_03250_),
    .B(_03251_),
    .Y(_03252_)
  );
  AOI22X1 _08746_ (
    .A( execution_unit_0.register_file_0.r1_5_ ),
    .B(_03113_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_5_ ),
    .Y(_02362_)
  );
  AOI22X1 _08747_ (
    .A( execution_unit_0.register_file_0.r4_5_ ),
    .B(_03126_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_5_ ),
    .Y(_02363_)
  );
  NAND2X1 _08748_ (
    .A(_02362_),
    .B(_02363_),
    .Y(_02364_)
  );
  NOR2X1 _08749_ (
    .A(_03252_),
    .B(_02364_),
    .Y(_02365_)
  );
  AOI22X1 _08750_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .B(_03117_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02366_)
  );
  AOI22X1 _08751_ (
    .A( execution_unit_0.register_file_0.r9_5_ ),
    .B(_03114_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_5_ ),
    .Y(_02367_)
  );
  NAND2X1 _08752_ (
    .A(_02366_),
    .B(_02367_),
    .Y(_02368_)
  );
  AOI22X1 _08753_ (
    .A( execution_unit_0.register_file_0.r11_5_ ),
    .B(_03112_),
    .C(_03115_),
    .D( execution_unit_0.register_file_0.r10_5_ ),
    .Y(_02369_)
  );
  AOI22X1 _08754_ (
    .A( execution_unit_0.register_file_0.r8_5_ ),
    .B(_03116_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02370_)
  );
  NAND2X1 _08755_ (
    .A(_02369_),
    .B(_02370_),
    .Y(_02371_)
  );
  NOR2X1 _08756_ (
    .A(_02368_),
    .B(_02371_),
    .Y(_02372_)
  );
  NAND2X1 _08757_ (
    .A(_02365_),
    .B(_02372_),
    .Y( execution_unit_0.reg_src_5_ )
  );
  INVX1 _08758_ (
    .A( execution_unit_0.reg_src_5_ ),
    .Y(_02373_)
  );
  AOI22X1 _08759_ (
    .A( dbg_0.UNUSED_pc_4_ ),
    .B(_03117_),
    .C(_03216_),
    .D( execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02374_)
  );
  AOI22X1 _08760_ (
    .A( execution_unit_0.register_file_0.r14_4_ ),
    .B(_03123_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02375_)
  );
  AOI22X1 _08761_ (
    .A( execution_unit_0.register_file_0.r1_4_ ),
    .B(_03113_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_4_ ),
    .Y(_02376_)
  );
  AOI22X1 _08762_ (
    .A( execution_unit_0.register_file_0.r10_4_ ),
    .B(_03115_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02377_)
  );
  AND2X1 _08763_ (
    .A(_02376_),
    .B(_02377_),
    .Y(_02378_)
  );
  NAND3X1 _08764_ (
    .A(_02374_),
    .B(_02375_),
    .C(_02378_),
    .Y(_02379_)
  );
  AOI22X1 _08765_ (
    .A( execution_unit_0.register_file_0.r13_4_ ),
    .B(_03111_),
    .C(_03114_),
    .D( execution_unit_0.register_file_0.r9_4_ ),
    .Y(_02380_)
  );
  AOI22X1 _08766_ (
    .A( execution_unit_0.register_file_0.r5_4_ ),
    .B(_03122_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_4_ ),
    .Y(_02381_)
  );
  AOI22X1 _08767_ (
    .A( execution_unit_0.register_file_0.r11_4_ ),
    .B(_03112_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_4_ ),
    .Y(_02382_)
  );
  AND2X1 _08768_ (
    .A(_02381_),
    .B(_02382_),
    .Y(_02383_)
  );
  AOI22X1 _08769_ (
    .A( execution_unit_0.register_file_0.r15_4_ ),
    .B(_03119_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_4_ ),
    .Y(_02384_)
  );
  NAND3X1 _08770_ (
    .A(_02380_),
    .B(_02383_),
    .C(_02384_),
    .Y(_02385_)
  );
  NOR2X1 _08771_ (
    .A(_02379_),
    .B(_02385_),
    .Y(_02386_)
  );
  INVX1 _08772_ (
    .A(_02386_),
    .Y( execution_unit_0.reg_src_4_ )
  );
  AOI22X1 _08773_ (
    .A( dbg_0.UNUSED_pc_3_ ),
    .B(_03117_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02387_)
  );
  AOI22X1 _08774_ (
    .A( execution_unit_0.register_file_0.r15_3_ ),
    .B(_03119_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_3_ ),
    .Y(_02388_)
  );
  AND2X1 _08775_ (
    .A(_02387_),
    .B(_02388_),
    .Y(_02389_)
  );
  AOI22X1 _08776_ (
    .A( execution_unit_0.register_file_0.r5_3_ ),
    .B(_03122_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_3_ ),
    .Y(_02390_)
  );
  AOI22X1 _08777_ (
    .A( execution_unit_0.register_file_0.r9_3_ ),
    .B(_03114_),
    .C(_03124_),
    .D( execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02391_)
  );
  NAND3X1 _08778_ (
    .A(_02389_),
    .B(_02390_),
    .C(_02391_),
    .Y(_02392_)
  );
  AOI22X1 _08779_ (
    .A( execution_unit_0.register_file_0.r11_3_ ),
    .B(_03112_),
    .C(_03216_),
    .D( execution_unit_0.gie ),
    .Y(_02393_)
  );
  AOI22X1 _08780_ (
    .A( execution_unit_0.register_file_0.r10_3_ ),
    .B(_03115_),
    .C(_03116_),
    .D( execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02394_)
  );
  AOI22X1 _08781_ (
    .A( execution_unit_0.register_file_0.r1_3_ ),
    .B(_03113_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_3_ ),
    .Y(_02395_)
  );
  AOI22X1 _08782_ (
    .A( execution_unit_0.register_file_0.r13_3_ ),
    .B(_03111_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_3_ ),
    .Y(_02396_)
  );
  AND2X1 _08783_ (
    .A(_02395_),
    .B(_02396_),
    .Y(_02397_)
  );
  NAND3X1 _08784_ (
    .A(_02393_),
    .B(_02394_),
    .C(_02397_),
    .Y(_02398_)
  );
  NOR2X1 _08785_ (
    .A(_02392_),
    .B(_02398_),
    .Y(_02399_)
  );
  INVX1 _08786_ (
    .A(_02399_),
    .Y( execution_unit_0.reg_src_3_ )
  );
  NAND2X1 _08787_ (
    .A( execution_unit_0.register_file_0.r10_2_ ),
    .B(_03115_),
    .Y(_02400_)
  );
  NAND2X1 _08788_ (
    .A( execution_unit_0.register_file_0.r11_2_ ),
    .B(_03112_),
    .Y(_02401_)
  );
  AOI22X1 _08789_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .B(_03117_),
    .C(_03122_),
    .D( execution_unit_0.register_file_0.r5_2_ ),
    .Y(_02402_)
  );
  AOI22X1 _08790_ (
    .A( execution_unit_0.register_file_0.r8_2_ ),
    .B(_03116_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_2_ ),
    .Y(_02403_)
  );
  NAND2X1 _08791_ (
    .A(_02400_),
    .B(_02403_),
    .Y(_02404_)
  );
  AOI22X1 _08792_ (
    .A( execution_unit_0.register_file_0.r6_2_ ),
    .B(_03124_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_2_ ),
    .Y(_02405_)
  );
  AOI22X1 _08793_ (
    .A( execution_unit_0.register_file_0.r9_2_ ),
    .B(_03114_),
    .C(_03125_),
    .D( execution_unit_0.register_file_0.r12_2_ ),
    .Y(_02406_)
  );
  AOI22X1 _08794_ (
    .A( execution_unit_0.register_file_0.r13_2_ ),
    .B(_03111_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_2_ ),
    .Y(_02407_)
  );
  NAND2X1 _08795_ (
    .A(_02406_),
    .B(_02407_),
    .Y(_02408_)
  );
  AOI22X1 _08796_ (
    .A( execution_unit_0.register_file_0.r1_2_ ),
    .B(_03113_),
    .C(_03216_),
    .D( execution_unit_0.alu_0.status_2_ ),
    .Y(_02409_)
  );
  NAND2X1 _08797_ (
    .A(_02401_),
    .B(_02409_),
    .Y(_02410_)
  );
  NOR2X1 _08798_ (
    .A(_02404_),
    .B(_02410_),
    .Y(_02411_)
  );
  AOI22X1 _08799_ (
    .A( execution_unit_0.register_file_0.r7_2_ ),
    .B(_03120_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_2_ ),
    .Y(_02412_)
  );
  NAND3X1 _08800_ (
    .A(_02402_),
    .B(_02405_),
    .C(_02412_),
    .Y(_02413_)
  );
  NOR2X1 _08801_ (
    .A(_02408_),
    .B(_02413_),
    .Y(_02414_)
  );
  AND2X1 _08802_ (
    .A(_02411_),
    .B(_02414_),
    .Y(_02415_)
  );
  INVX1 _08803_ (
    .A(_02415_),
    .Y( execution_unit_0.reg_src_2_ )
  );
  NAND3X1 _08804_ (
    .A( execution_unit_0.register_file_0.r6_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_6_ ),
    .Y(_02416_)
  );
  OAI21X1 _08805_ (
    .A(_03103_),
    .B(_03127_),
    .C(_02416_),
    .Y(_02417_)
  );
  OAI21X1 _08806_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .C( execution_unit_0.alu_0.status_1_ ),
    .Y(_02418_)
  );
  NAND3X1 _08807_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_0_ ),
    .C( dbg_0.UNUSED_pc_1_ ),
    .Y(_02419_)
  );
  AOI22X1 _08808_ (
    .A( execution_unit_0.register_file_0.r10_1_ ),
    .B(_03115_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02420_)
  );
  NAND2X1 _08809_ (
    .A( execution_unit_0.register_file_0.r11_1_ ),
    .B(_03112_),
    .Y(_02421_)
  );
  NAND3X1 _08810_ (
    .A( execution_unit_0.register_file_0.r12_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_12_ ),
    .Y(_02422_)
  );
  NAND3X1 _08811_ (
    .A( execution_unit_0.register_file_0.r15_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_15_ ),
    .Y(_02423_)
  );
  NAND3X1 _08812_ (
    .A( execution_unit_0.register_file_0.r8_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_8_ ),
    .Y(_02424_)
  );
  NAND3X1 _08813_ (
    .A( execution_unit_0.register_file_0.r5_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_5_ ),
    .Y(_02425_)
  );
  NAND3X1 _08814_ (
    .A( execution_unit_0.register_file_0.r9_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_9_ ),
    .Y(_02426_)
  );
  NAND3X1 _08815_ (
    .A( execution_unit_0.register_file_0.r3_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_3_ ),
    .Y(_02427_)
  );
  NAND3X1 _08816_ (
    .A( execution_unit_0.register_file_0.r13_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_13_ ),
    .Y(_02428_)
  );
  NAND3X1 _08817_ (
    .A( execution_unit_0.register_file_0.r1_1_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_1_ ),
    .Y(_02429_)
  );
  AND2X1 _08818_ (
    .A( execution_unit_0.register_file_0.r14_1_ ),
    .B(_03123_),
    .Y(_02430_)
  );
  NAND3X1 _08819_ (
    .A(_02419_),
    .B(_02423_),
    .C(_02429_),
    .Y(_02431_)
  );
  NAND3X1 _08820_ (
    .A(_02418_),
    .B(_02425_),
    .C(_02427_),
    .Y(_02432_)
  );
  NOR3X1 _08821_ (
    .A(_02417_),
    .B(_02431_),
    .C(_02432_),
    .Y(_02433_)
  );
  NAND2X1 _08822_ (
    .A(_02426_),
    .B(_02428_),
    .Y(_02434_)
  );
  NAND2X1 _08823_ (
    .A(_02422_),
    .B(_02424_),
    .Y(_02435_)
  );
  NOR3X1 _08824_ (
    .A(_02430_),
    .B(_02434_),
    .C(_02435_),
    .Y(_02436_)
  );
  AND2X1 _08825_ (
    .A(_02420_),
    .B(_02421_),
    .Y(_02437_)
  );
  AND2X1 _08826_ (
    .A(_02436_),
    .B(_02437_),
    .Y(_02438_)
  );
  NAND3X1 _08827_ (
    .A(_02433_),
    .B(_02436_),
    .C(_02437_),
    .Y( execution_unit_0.reg_src_1_ )
  );
  OAI21X1 _08828_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_03106_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_02439_)
  );
  INVX1 _08829_ (
    .A(_02439_),
    .Y(_02440_)
  );
  NAND2X1 _08830_ (
    .A( execution_unit_0.register_file_0.r9_0_ ),
    .B(_03114_),
    .Y(_02441_)
  );
  NAND2X1 _08831_ (
    .A( execution_unit_0.register_file_0.r11_0_ ),
    .B(_03112_),
    .Y(_02442_)
  );
  NAND2X1 _08832_ (
    .A( execution_unit_0.register_file_0.r14_0_ ),
    .B(_03123_),
    .Y(_02443_)
  );
  AOI22X1 _08833_ (
    .A( execution_unit_0.register_file_0.r13_0_ ),
    .B(_03111_),
    .C(_03119_),
    .D( execution_unit_0.register_file_0.r15_0_ ),
    .Y(_02444_)
  );
  AOI22X1 _08834_ (
    .A( execution_unit_0.register_file_0.r6_0_ ),
    .B(_03124_),
    .C(_03216_),
    .D( execution_unit_0.alu_0.status_0_ ),
    .Y(_02445_)
  );
  NAND3X1 _08835_ (
    .A(_03105_),
    .B( execution_unit_0.inst_src_0_ ),
    .C( dbg_0.UNUSED_pc_0_ ),
    .Y(_02446_)
  );
  NAND3X1 _08836_ (
    .A( execution_unit_0.register_file_0.r12_0_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_12_ ),
    .Y(_02447_)
  );
  NAND3X1 _08837_ (
    .A( execution_unit_0.register_file_0.r8_0_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_8_ ),
    .Y(_02448_)
  );
  NAND3X1 _08838_ (
    .A( execution_unit_0.register_file_0.r5_0_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_5_ ),
    .Y(_02449_)
  );
  NAND3X1 _08839_ (
    .A( execution_unit_0.register_file_0.r10_0_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_10_ ),
    .Y(_02450_)
  );
  NAND3X1 _08840_ (
    .A( execution_unit_0.register_file_0.r3_0_ ),
    .B(_03105_),
    .C( execution_unit_0.inst_src_3_ ),
    .Y(_02451_)
  );
  AOI22X1 _08841_ (
    .A( execution_unit_0.register_file_0.r7_0_ ),
    .B(_03120_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_0_ ),
    .Y(_02452_)
  );
  AND2X1 _08842_ (
    .A(_02447_),
    .B(_02450_),
    .Y(_02453_)
  );
  NAND3X1 _08843_ (
    .A(_02441_),
    .B(_02444_),
    .C(_02453_),
    .Y(_02454_)
  );
  NAND3X1 _08844_ (
    .A(_02442_),
    .B(_02443_),
    .C(_02452_),
    .Y(_02455_)
  );
  AND2X1 _08845_ (
    .A(_02448_),
    .B(_02451_),
    .Y(_02456_)
  );
  AND2X1 _08846_ (
    .A(_02446_),
    .B(_02449_),
    .Y(_02457_)
  );
  NAND3X1 _08847_ (
    .A(_02445_),
    .B(_02456_),
    .C(_02457_),
    .Y(_02458_)
  );
  NOR3X1 _08848_ (
    .A(_02454_),
    .B(_02455_),
    .C(_02458_),
    .Y(_02459_)
  );
  INVX1 _08849_ (
    .A(_02459_),
    .Y( execution_unit_0.reg_src_0_ )
  );
  NAND2X1 _08850_ (
    .A(_02440_),
    .B(_02459_),
    .Y(_02460_)
  );
  AOI22X1 _08851_ (
    .A(_02433_),
    .B(_02438_),
    .C(_02440_),
    .D(_02459_),
    .Y(_02461_)
  );
  OAI21X1 _08852_ (
    .A(_02439_),
    .B( execution_unit_0.reg_src_0_ ),
    .C( execution_unit_0.reg_src_1_ ),
    .Y(_02462_)
  );
  NOR3X1 _08853_ (
    .A(_02399_),
    .B(_02415_),
    .C(_02462_),
    .Y(_02463_)
  );
  NAND3X1 _08854_ (
    .A( execution_unit_0.reg_src_3_ ),
    .B( execution_unit_0.reg_src_2_ ),
    .C(_02461_),
    .Y(_02464_)
  );
  NOR3X1 _08855_ (
    .A(_02373_),
    .B(_02386_),
    .C(_02464_),
    .Y(_02465_)
  );
  NAND3X1 _08856_ (
    .A( execution_unit_0.reg_src_5_ ),
    .B( execution_unit_0.reg_src_4_ ),
    .C(_02463_),
    .Y(_02466_)
  );
  NOR3X1 _08857_ (
    .A(_03236_),
    .B(_03249_),
    .C(_02466_),
    .Y(_02467_)
  );
  NAND3X1 _08858_ (
    .A( execution_unit_0.reg_src_7_ ),
    .B( execution_unit_0.reg_src_6_ ),
    .C(_02465_),
    .Y(_02468_)
  );
  NOR3X1 _08859_ (
    .A(_03209_),
    .B(_03223_),
    .C(_02468_),
    .Y(_02469_)
  );
  NAND3X1 _08860_ (
    .A( execution_unit_0.reg_src_9_ ),
    .B( execution_unit_0.reg_src_8_ ),
    .C(_02467_),
    .Y(_02470_)
  );
  NOR3X1 _08861_ (
    .A(_03182_),
    .B(_03195_),
    .C(_02470_),
    .Y(_02471_)
  );
  NAND3X1 _08862_ (
    .A( execution_unit_0.reg_src_11_ ),
    .B( execution_unit_0.reg_src_10_ ),
    .C(_02469_),
    .Y(_02472_)
  );
  NOR3X1 _08863_ (
    .A(_03153_),
    .B(_03168_),
    .C(_02472_),
    .Y(_02473_)
  );
  NAND3X1 _08864_ (
    .A( execution_unit_0.reg_src_13_ ),
    .B( execution_unit_0.reg_src_12_ ),
    .C(_02471_),
    .Y(_02474_)
  );
  NAND2X1 _08865_ (
    .A( execution_unit_0.register_file_0.r12_15_ ),
    .B(_03125_),
    .Y(_02475_)
  );
  NAND2X1 _08866_ (
    .A( execution_unit_0.register_file_0.r8_15_ ),
    .B(_03116_),
    .Y(_02476_)
  );
  AOI22X1 _08867_ (
    .A( execution_unit_0.register_file_0.r6_15_ ),
    .B(_03124_),
    .C(_03128_),
    .D( execution_unit_0.register_file_0.r3_15_ ),
    .Y(_02477_)
  );
  AOI22X1 _08868_ (
    .A( execution_unit_0.register_file_0.r9_15_ ),
    .B(_03114_),
    .C(_03120_),
    .D( execution_unit_0.register_file_0.r7_15_ ),
    .Y(_02478_)
  );
  AOI22X1 _08869_ (
    .A( execution_unit_0.register_file_0.r1_15_ ),
    .B(_03113_),
    .C(_03117_),
    .D( dbg_0.UNUSED_pc_15_ ),
    .Y(_02479_)
  );
  AOI22X1 _08870_ (
    .A( execution_unit_0.register_file_0.r15_15_ ),
    .B(_03119_),
    .C(_03123_),
    .D( execution_unit_0.register_file_0.r14_15_ ),
    .Y(_02480_)
  );
  AOI22X1 _08871_ (
    .A( execution_unit_0.register_file_0.r13_15_ ),
    .B(_03111_),
    .C(_03115_),
    .D( execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02481_)
  );
  NAND2X1 _08872_ (
    .A(_02480_),
    .B(_02481_),
    .Y(_02482_)
  );
  AOI21X1 _08873_ (
    .A( execution_unit_0.register_file_0.r11_15_ ),
    .B(_03112_),
    .C(_02482_),
    .Y(_02483_)
  );
  NAND3X1 _08874_ (
    .A(_02475_),
    .B(_02476_),
    .C(_02479_),
    .Y(_02484_)
  );
  AOI22X1 _08875_ (
    .A( execution_unit_0.register_file_0.r5_15_ ),
    .B(_03122_),
    .C(_03126_),
    .D( execution_unit_0.register_file_0.r4_15_ ),
    .Y(_02485_)
  );
  NAND3X1 _08876_ (
    .A(_02477_),
    .B(_02478_),
    .C(_02485_),
    .Y(_02486_)
  );
  NOR2X1 _08877_ (
    .A(_02484_),
    .B(_02486_),
    .Y(_02487_)
  );
  NAND2X1 _08878_ (
    .A(_02483_),
    .B(_02487_),
    .Y( execution_unit_0.reg_src_15_ )
  );
  INVX1 _08879_ (
    .A( execution_unit_0.reg_src_15_ ),
    .Y(_02488_)
  );
  NAND3X1 _08880_ (
    .A( execution_unit_0.reg_src_14_ ),
    .B(_02473_),
    .C( execution_unit_0.reg_src_15_ ),
    .Y(_02489_)
  );
  OAI21X1 _08881_ (
    .A(_03140_),
    .B(_02474_),
    .C(_02488_),
    .Y(_02490_)
  );
  NAND2X1 _08882_ (
    .A(_02489_),
    .B(_02490_),
    .Y(_02491_)
  );
  AOI21X1 _08883_ (
    .A(_02489_),
    .B(_02490_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02492_)
  );
  AOI21X1 _08884_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03113_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02493_)
  );
  AND2X1 _08885_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.reg_dest_wr ),
    .Y(_02494_)
  );
  NAND2X1 _08886_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.reg_dest_wr ),
    .Y(_02495_)
  );
  NOR2X1 _08887_ (
    .A(_02493_),
    .B(_02494_),
    .Y(_02496_)
  );
  OAI21X1 _08888_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_15_ ),
    .C(_02496_),
    .Y(_02497_)
  );
  AND2X1 _08889_ (
    .A(_02493_),
    .B(_02495_),
    .Y(_02498_)
  );
  AND2X1 _08890_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .Y( execution_unit_0.pc_sw_15_ )
  );
  INVX1 _08891_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .Y(_02499_)
  );
  AOI22X1 _08892_ (
    .A( execution_unit_0.register_file_0.r1_15_ ),
    .B(_02498_),
    .C( execution_unit_0.pc_sw_15_ ),
    .D(_02494_),
    .Y(_02500_)
  );
  OAI21X1 _08893_ (
    .A(_02492_),
    .B(_02497_),
    .C(_02500_),
    .Y(_02361_)
  );
  XNOR2X1 _08894_ (
    .A(_03140_),
    .B(_02473_),
    .Y(_02501_)
  );
  NOR2X1 _08895_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02501_),
    .Y(_02502_)
  );
  OAI21X1 _08896_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .C(_02496_),
    .Y(_02503_)
  );
  AND2X1 _08897_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .Y( execution_unit_0.pc_sw_14_ )
  );
  INVX1 _08898_ (
    .A( execution_unit_0.pc_sw_14_ ),
    .Y(_02504_)
  );
  AOI22X1 _08899_ (
    .A( execution_unit_0.register_file_0.r1_14_ ),
    .B(_02498_),
    .C( execution_unit_0.pc_sw_14_ ),
    .D(_02494_),
    .Y(_02505_)
  );
  OAI21X1 _08900_ (
    .A(_02502_),
    .B(_02503_),
    .C(_02505_),
    .Y(_02360_)
  );
  OAI21X1 _08901_ (
    .A(_03168_),
    .B(_02472_),
    .C(_03153_),
    .Y(_02506_)
  );
  NAND2X1 _08902_ (
    .A(_02474_),
    .B(_02506_),
    .Y(_02507_)
  );
  AOI21X1 _08903_ (
    .A(_02474_),
    .B(_02506_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02508_)
  );
  OAI21X1 _08904_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .C(_02496_),
    .Y(_02509_)
  );
  AND2X1 _08905_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_13_ ),
    .Y( execution_unit_0.pc_sw_13_ )
  );
  INVX1 _08906_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .Y(_02510_)
  );
  AOI22X1 _08907_ (
    .A( execution_unit_0.register_file_0.r1_13_ ),
    .B(_02498_),
    .C( execution_unit_0.pc_sw_13_ ),
    .D(_02494_),
    .Y(_02511_)
  );
  OAI21X1 _08908_ (
    .A(_02508_),
    .B(_02509_),
    .C(_02511_),
    .Y(_02359_)
  );
  XNOR2X1 _08909_ (
    .A( execution_unit_0.reg_src_12_ ),
    .B(_02471_),
    .Y(_02512_)
  );
  OAI21X1 _08910_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_12_ ),
    .C(_02496_),
    .Y(_02513_)
  );
  AOI21X1 _08911_ (
    .A(_03104_),
    .B(_02512_),
    .C(_02513_),
    .Y(_02514_)
  );
  NAND2X1 _08912_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_12_ ),
    .Y(_02515_)
  );
  INVX1 _08913_ (
    .A(_02515_),
    .Y( execution_unit_0.pc_sw_12_ )
  );
  AOI21X1 _08914_ (
    .A( execution_unit_0.register_file_0.r1_12_ ),
    .B(_02498_),
    .C(_02514_),
    .Y(_02516_)
  );
  OAI21X1 _08915_ (
    .A(_02495_),
    .B(_02515_),
    .C(_02516_),
    .Y(_02358_)
  );
  OAI21X1 _08916_ (
    .A(_03195_),
    .B(_02470_),
    .C(_03182_),
    .Y(_02517_)
  );
  NAND2X1 _08917_ (
    .A(_02472_),
    .B(_02517_),
    .Y(_02518_)
  );
  OAI21X1 _08918_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .C(_02496_),
    .Y(_02519_)
  );
  AOI21X1 _08919_ (
    .A(_03104_),
    .B(_02518_),
    .C(_02519_),
    .Y(_02520_)
  );
  AND2X1 _08920_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_11_ ),
    .Y( execution_unit_0.pc_sw_11_ )
  );
  INVX1 _08921_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .Y(_02521_)
  );
  AOI21X1 _08922_ (
    .A( execution_unit_0.register_file_0.r1_11_ ),
    .B(_02498_),
    .C(_02520_),
    .Y(_02522_)
  );
  OAI21X1 _08923_ (
    .A(_02495_),
    .B(_02521_),
    .C(_02522_),
    .Y(_02357_)
  );
  XNOR2X1 _08924_ (
    .A(_03195_),
    .B(_02469_),
    .Y(_02523_)
  );
  NOR2X1 _08925_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02523_),
    .Y(_02524_)
  );
  OAI21X1 _08926_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_10_ ),
    .C(_02496_),
    .Y(_02525_)
  );
  AND2X1 _08927_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_10_ ),
    .Y( execution_unit_0.pc_sw_10_ )
  );
  INVX1 _08928_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .Y(_02526_)
  );
  AOI22X1 _08929_ (
    .A( execution_unit_0.register_file_0.r1_10_ ),
    .B(_02498_),
    .C( execution_unit_0.pc_sw_10_ ),
    .D(_02494_),
    .Y(_02527_)
  );
  OAI21X1 _08930_ (
    .A(_02524_),
    .B(_02525_),
    .C(_02527_),
    .Y(_02356_)
  );
  OAI21X1 _08931_ (
    .A(_03223_),
    .B(_02468_),
    .C(_03209_),
    .Y(_02528_)
  );
  NAND2X1 _08932_ (
    .A(_02470_),
    .B(_02528_),
    .Y(_02529_)
  );
  OAI21X1 _08933_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_9_ ),
    .C(_02496_),
    .Y(_02530_)
  );
  AOI21X1 _08934_ (
    .A(_03104_),
    .B(_02529_),
    .C(_02530_),
    .Y(_02531_)
  );
  AND2X1 _08935_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_9_ ),
    .Y( execution_unit_0.pc_sw_9_ )
  );
  INVX1 _08936_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .Y(_02532_)
  );
  AOI21X1 _08937_ (
    .A( execution_unit_0.register_file_0.r1_9_ ),
    .B(_02498_),
    .C(_02531_),
    .Y(_02533_)
  );
  OAI21X1 _08938_ (
    .A(_02495_),
    .B(_02532_),
    .C(_02533_),
    .Y(_02355_)
  );
  XNOR2X1 _08939_ (
    .A(_03223_),
    .B(_02467_),
    .Y(_02534_)
  );
  NOR2X1 _08940_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02534_),
    .Y(_02535_)
  );
  OAI21X1 _08941_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_8_ ),
    .C(_02496_),
    .Y(_02536_)
  );
  NAND2X1 _08942_ (
    .A(_03108_),
    .B( execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_02537_)
  );
  INVX1 _08943_ (
    .A(_02537_),
    .Y( execution_unit_0.pc_sw_8_ )
  );
  AOI22X1 _08944_ (
    .A( execution_unit_0.register_file_0.r1_8_ ),
    .B(_02498_),
    .C( execution_unit_0.pc_sw_8_ ),
    .D(_02494_),
    .Y(_02538_)
  );
  OAI21X1 _08945_ (
    .A(_02535_),
    .B(_02536_),
    .C(_02538_),
    .Y(_02354_)
  );
  OAI21X1 _08946_ (
    .A(_03249_),
    .B(_02466_),
    .C(_03236_),
    .Y(_02539_)
  );
  NAND2X1 _08947_ (
    .A(_02468_),
    .B(_02539_),
    .Y(_02540_)
  );
  OAI21X1 _08948_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .C(_02496_),
    .Y(_02541_)
  );
  AOI21X1 _08949_ (
    .A(_03104_),
    .B(_02540_),
    .C(_02541_),
    .Y(_02542_)
  );
  AOI21X1 _08950_ (
    .A( execution_unit_0.register_file_0.r1_7_ ),
    .B(_02498_),
    .C(_02542_),
    .Y(_02543_)
  );
  OAI21X1 _08951_ (
    .A(_03094_),
    .B(_02495_),
    .C(_02543_),
    .Y(_02353_)
  );
  XNOR2X1 _08952_ (
    .A( execution_unit_0.reg_src_6_ ),
    .B(_02465_),
    .Y(_02544_)
  );
  OAI21X1 _08953_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_6_ ),
    .C(_02496_),
    .Y(_02545_)
  );
  AOI21X1 _08954_ (
    .A(_03104_),
    .B(_02544_),
    .C(_02545_),
    .Y(_02546_)
  );
  AOI21X1 _08955_ (
    .A( execution_unit_0.register_file_0.r1_6_ ),
    .B(_02498_),
    .C(_02546_),
    .Y(_02547_)
  );
  OAI21X1 _08956_ (
    .A(_03095_),
    .B(_02495_),
    .C(_02547_),
    .Y(_02352_)
  );
  OAI21X1 _08957_ (
    .A(_02386_),
    .B(_02464_),
    .C(_02373_),
    .Y(_02548_)
  );
  NAND2X1 _08958_ (
    .A(_02466_),
    .B(_02548_),
    .Y(_02549_)
  );
  OAI21X1 _08959_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_5_ ),
    .C(_02496_),
    .Y(_02550_)
  );
  AOI21X1 _08960_ (
    .A(_03104_),
    .B(_02549_),
    .C(_02550_),
    .Y(_02551_)
  );
  AOI21X1 _08961_ (
    .A( execution_unit_0.register_file_0.r1_5_ ),
    .B(_02498_),
    .C(_02551_),
    .Y(_02552_)
  );
  OAI21X1 _08962_ (
    .A(_03096_),
    .B(_02495_),
    .C(_02552_),
    .Y(_02351_)
  );
  XNOR2X1 _08963_ (
    .A( execution_unit_0.reg_src_4_ ),
    .B(_02463_),
    .Y(_02553_)
  );
  OAI21X1 _08964_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .C(_02496_),
    .Y(_02554_)
  );
  AOI21X1 _08965_ (
    .A(_03104_),
    .B(_02553_),
    .C(_02554_),
    .Y(_02555_)
  );
  AOI21X1 _08966_ (
    .A( execution_unit_0.register_file_0.r1_4_ ),
    .B(_02498_),
    .C(_02555_),
    .Y(_02556_)
  );
  OAI21X1 _08967_ (
    .A(_03097_),
    .B(_02495_),
    .C(_02556_),
    .Y(_02350_)
  );
  OAI21X1 _08968_ (
    .A(_02415_),
    .B(_02462_),
    .C(_02399_),
    .Y(_02557_)
  );
  NAND2X1 _08969_ (
    .A(_02464_),
    .B(_02557_),
    .Y(_02558_)
  );
  OAI21X1 _08970_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_3_ ),
    .C(_02496_),
    .Y(_02559_)
  );
  AOI21X1 _08971_ (
    .A(_03104_),
    .B(_02558_),
    .C(_02559_),
    .Y(_02560_)
  );
  AOI21X1 _08972_ (
    .A( execution_unit_0.register_file_0.r1_3_ ),
    .B(_02498_),
    .C(_02560_),
    .Y(_02561_)
  );
  OAI21X1 _08973_ (
    .A(_03098_),
    .B(_02495_),
    .C(_02561_),
    .Y(_02349_)
  );
  XNOR2X1 _08974_ (
    .A(_02415_),
    .B(_02461_),
    .Y(_02562_)
  );
  NOR2X1 _08975_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02562_),
    .Y(_02563_)
  );
  OAI21X1 _08976_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .C(_02496_),
    .Y(_02564_)
  );
  AOI22X1 _08977_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02494_),
    .C(_02498_),
    .D( execution_unit_0.register_file_0.r1_2_ ),
    .Y(_02565_)
  );
  OAI21X1 _08978_ (
    .A(_02563_),
    .B(_02564_),
    .C(_02565_),
    .Y(_02348_)
  );
  XNOR2X1 _08979_ (
    .A( execution_unit_0.reg_src_1_ ),
    .B(_02460_),
    .Y(_02566_)
  );
  AND2X1 _08980_ (
    .A(_03104_),
    .B(_02566_),
    .Y(_02567_)
  );
  OAI21X1 _08981_ (
    .A(_03104_),
    .B( dbg_0.UNUSED_eu_mab_1_ ),
    .C(_02496_),
    .Y(_02568_)
  );
  AOI22X1 _08982_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02494_),
    .C(_02498_),
    .D( execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02569_)
  );
  OAI21X1 _08983_ (
    .A(_02567_),
    .B(_02568_),
    .C(_02569_),
    .Y(_02347_)
  );
  AOI21X1 _08984_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.reg_sr_wr ),
    .Y(_02570_)
  );
  MUX2X1 _08985_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.alu_0.alu_out_0_ ),
    .S(_02570_),
    .Y(_02571_)
  );
  OAI21X1 _08986_ (
    .A(_03107_),
    .B( execution_unit_0.alu_0.alu_stat_0_ ),
    .C(_03105_),
    .Y(_02572_)
  );
  AOI21X1 _08987_ (
    .A(_03107_),
    .B(_02571_),
    .C(_02572_),
    .Y(_02346_)
  );
  NAND2X1 _08988_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_3_ ),
    .Y(_02573_)
  );
  NAND2X1 _08989_ (
    .A( execution_unit_0.register_file_0.r3_15_ ),
    .B(_02573_),
    .Y(_02574_)
  );
  OAI21X1 _08990_ (
    .A(_02499_),
    .B(_02573_),
    .C(_02574_),
    .Y(_02345_)
  );
  NAND2X1 _08991_ (
    .A( execution_unit_0.register_file_0.r3_14_ ),
    .B(_02573_),
    .Y(_02575_)
  );
  OAI21X1 _08992_ (
    .A(_02504_),
    .B(_02573_),
    .C(_02575_),
    .Y(_02344_)
  );
  NAND2X1 _08993_ (
    .A( execution_unit_0.register_file_0.r3_13_ ),
    .B(_02573_),
    .Y(_02576_)
  );
  OAI21X1 _08994_ (
    .A(_02510_),
    .B(_02573_),
    .C(_02576_),
    .Y(_02343_)
  );
  NAND2X1 _08995_ (
    .A( execution_unit_0.register_file_0.r3_12_ ),
    .B(_02573_),
    .Y(_02577_)
  );
  OAI21X1 _08996_ (
    .A(_02515_),
    .B(_02573_),
    .C(_02577_),
    .Y(_02342_)
  );
  NAND2X1 _08997_ (
    .A( execution_unit_0.register_file_0.r3_11_ ),
    .B(_02573_),
    .Y(_02578_)
  );
  OAI21X1 _08998_ (
    .A(_02521_),
    .B(_02573_),
    .C(_02578_),
    .Y(_02341_)
  );
  NAND2X1 _08999_ (
    .A( execution_unit_0.register_file_0.r3_10_ ),
    .B(_02573_),
    .Y(_02579_)
  );
  OAI21X1 _09000_ (
    .A(_02526_),
    .B(_02573_),
    .C(_02579_),
    .Y(_02340_)
  );
  NAND2X1 _09001_ (
    .A( execution_unit_0.register_file_0.r3_9_ ),
    .B(_02573_),
    .Y(_02580_)
  );
  OAI21X1 _09002_ (
    .A(_02532_),
    .B(_02573_),
    .C(_02580_),
    .Y(_02339_)
  );
  NAND2X1 _09003_ (
    .A( execution_unit_0.register_file_0.r3_8_ ),
    .B(_02573_),
    .Y(_02581_)
  );
  OAI21X1 _09004_ (
    .A(_02537_),
    .B(_02573_),
    .C(_02581_),
    .Y(_02338_)
  );
  NAND2X1 _09005_ (
    .A( execution_unit_0.register_file_0.r3_7_ ),
    .B(_02573_),
    .Y(_02582_)
  );
  OAI21X1 _09006_ (
    .A(_03094_),
    .B(_02573_),
    .C(_02582_),
    .Y(_02337_)
  );
  NAND2X1 _09007_ (
    .A( execution_unit_0.register_file_0.r3_6_ ),
    .B(_02573_),
    .Y(_02583_)
  );
  OAI21X1 _09008_ (
    .A(_03095_),
    .B(_02573_),
    .C(_02583_),
    .Y(_02336_)
  );
  NAND2X1 _09009_ (
    .A( execution_unit_0.register_file_0.r3_5_ ),
    .B(_02573_),
    .Y(_02584_)
  );
  OAI21X1 _09010_ (
    .A(_03096_),
    .B(_02573_),
    .C(_02584_),
    .Y(_02335_)
  );
  NAND2X1 _09011_ (
    .A( execution_unit_0.register_file_0.r3_4_ ),
    .B(_02573_),
    .Y(_02585_)
  );
  OAI21X1 _09012_ (
    .A(_03097_),
    .B(_02573_),
    .C(_02585_),
    .Y(_02334_)
  );
  NAND2X1 _09013_ (
    .A( execution_unit_0.register_file_0.r3_3_ ),
    .B(_02573_),
    .Y(_02586_)
  );
  OAI21X1 _09014_ (
    .A(_03098_),
    .B(_02573_),
    .C(_02586_),
    .Y(_02333_)
  );
  NAND2X1 _09015_ (
    .A( execution_unit_0.register_file_0.r3_2_ ),
    .B(_02573_),
    .Y(_02587_)
  );
  OAI21X1 _09016_ (
    .A(_03099_),
    .B(_02573_),
    .C(_02587_),
    .Y(_02332_)
  );
  NAND2X1 _09017_ (
    .A( execution_unit_0.register_file_0.r3_1_ ),
    .B(_02573_),
    .Y(_02588_)
  );
  OAI21X1 _09018_ (
    .A(_03100_),
    .B(_02573_),
    .C(_02588_),
    .Y(_02331_)
  );
  NAND2X1 _09019_ (
    .A( execution_unit_0.register_file_0.r3_0_ ),
    .B(_02573_),
    .Y(_02589_)
  );
  OAI21X1 _09020_ (
    .A(_03101_),
    .B(_02573_),
    .C(_02589_),
    .Y(_02330_)
  );
  AND2X1 _09021_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_4_ ),
    .Y(_02590_)
  );
  NAND2X1 _09022_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_4_ ),
    .Y(_02591_)
  );
  NAND2X1 _09023_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03126_),
    .Y(_02592_)
  );
  NOR2X1 _09024_ (
    .A(_02590_),
    .B(_02592_),
    .Y(_02593_)
  );
  OR2X1 _09025_ (
    .A(_02590_),
    .B(_02592_),
    .Y(_02594_)
  );
  AOI21X1 _09026_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03126_),
    .C(_02590_),
    .Y(_02595_)
  );
  AOI22X1 _09027_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_15_ ),
    .Y(_02596_)
  );
  OAI21X1 _09028_ (
    .A(_02491_),
    .B(_02594_),
    .C(_02596_),
    .Y(_02329_)
  );
  AOI22X1 _09029_ (
    .A(_02501_),
    .B(_02593_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_14_ ),
    .Y(_02597_)
  );
  OAI21X1 _09030_ (
    .A(_02504_),
    .B(_02591_),
    .C(_02597_),
    .Y(_02328_)
  );
  AOI22X1 _09031_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_13_ ),
    .Y(_02598_)
  );
  OAI21X1 _09032_ (
    .A(_02507_),
    .B(_02594_),
    .C(_02598_),
    .Y(_02327_)
  );
  AOI22X1 _09033_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_12_ ),
    .Y(_02599_)
  );
  OAI21X1 _09034_ (
    .A(_02512_),
    .B(_02594_),
    .C(_02599_),
    .Y(_02326_)
  );
  AOI22X1 _09035_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_11_ ),
    .Y(_02600_)
  );
  OAI21X1 _09036_ (
    .A(_02518_),
    .B(_02594_),
    .C(_02600_),
    .Y(_02325_)
  );
  AOI22X1 _09037_ (
    .A(_02523_),
    .B(_02593_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_10_ ),
    .Y(_02601_)
  );
  OAI21X1 _09038_ (
    .A(_02526_),
    .B(_02591_),
    .C(_02601_),
    .Y(_02324_)
  );
  AOI22X1 _09039_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_9_ ),
    .Y(_02602_)
  );
  OAI21X1 _09040_ (
    .A(_02529_),
    .B(_02594_),
    .C(_02602_),
    .Y(_02323_)
  );
  AOI22X1 _09041_ (
    .A(_02534_),
    .B(_02593_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_8_ ),
    .Y(_02603_)
  );
  OAI21X1 _09042_ (
    .A(_02537_),
    .B(_02591_),
    .C(_02603_),
    .Y(_02322_)
  );
  AOI22X1 _09043_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_7_ ),
    .Y(_02604_)
  );
  OAI21X1 _09044_ (
    .A(_02540_),
    .B(_02594_),
    .C(_02604_),
    .Y(_02321_)
  );
  AOI22X1 _09045_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_6_ ),
    .Y(_02605_)
  );
  OAI21X1 _09046_ (
    .A(_02544_),
    .B(_02594_),
    .C(_02605_),
    .Y(_02320_)
  );
  AOI22X1 _09047_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_5_ ),
    .Y(_02606_)
  );
  OAI21X1 _09048_ (
    .A(_02549_),
    .B(_02594_),
    .C(_02606_),
    .Y(_02319_)
  );
  AOI22X1 _09049_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02607_)
  );
  OAI21X1 _09050_ (
    .A(_02553_),
    .B(_02594_),
    .C(_02607_),
    .Y(_02318_)
  );
  AOI22X1 _09051_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_3_ ),
    .Y(_02608_)
  );
  OAI21X1 _09052_ (
    .A(_02558_),
    .B(_02594_),
    .C(_02608_),
    .Y(_02317_)
  );
  NAND2X1 _09053_ (
    .A( execution_unit_0.register_file_0.r4_2_ ),
    .B(_02595_),
    .Y(_02609_)
  );
  AOI22X1 _09054_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02590_),
    .C(_02593_),
    .D(_02562_),
    .Y(_02610_)
  );
  NAND2X1 _09055_ (
    .A(_02609_),
    .B(_02610_),
    .Y(_02316_)
  );
  AOI22X1 _09056_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02590_),
    .C(_02595_),
    .D( execution_unit_0.register_file_0.r4_1_ ),
    .Y(_02611_)
  );
  OAI21X1 _09057_ (
    .A(_02566_),
    .B(_02594_),
    .C(_02611_),
    .Y(_02315_)
  );
  OAI21X1 _09058_ (
    .A(_03108_),
    .B(_03113_),
    .C( execution_unit_0.reg_src_0_ ),
    .Y(_02612_)
  );
  NAND2X1 _09059_ (
    .A(_02460_),
    .B(_02612_),
    .Y(_02613_)
  );
  NAND2X1 _09060_ (
    .A( execution_unit_0.register_file_0.r4_0_ ),
    .B(_02595_),
    .Y(_02614_)
  );
  AOI22X1 _09061_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02590_),
    .C(_02593_),
    .D(_02613_),
    .Y(_02615_)
  );
  NAND2X1 _09062_ (
    .A(_02614_),
    .B(_02615_),
    .Y(_02314_)
  );
  AND2X1 _09063_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_5_ ),
    .Y(_02616_)
  );
  NAND2X1 _09064_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_5_ ),
    .Y(_02617_)
  );
  NAND2X1 _09065_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03122_),
    .Y(_02618_)
  );
  NOR2X1 _09066_ (
    .A(_02616_),
    .B(_02618_),
    .Y(_02619_)
  );
  OR2X1 _09067_ (
    .A(_02616_),
    .B(_02618_),
    .Y(_02620_)
  );
  AOI21X1 _09068_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03122_),
    .C(_02616_),
    .Y(_02621_)
  );
  AOI22X1 _09069_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_15_ ),
    .Y(_02622_)
  );
  OAI21X1 _09070_ (
    .A(_02491_),
    .B(_02620_),
    .C(_02622_),
    .Y(_02313_)
  );
  AOI22X1 _09071_ (
    .A(_02501_),
    .B(_02619_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_14_ ),
    .Y(_02623_)
  );
  OAI21X1 _09072_ (
    .A(_02504_),
    .B(_02617_),
    .C(_02623_),
    .Y(_02312_)
  );
  AOI22X1 _09073_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_13_ ),
    .Y(_02624_)
  );
  OAI21X1 _09074_ (
    .A(_02507_),
    .B(_02620_),
    .C(_02624_),
    .Y(_02311_)
  );
  AOI22X1 _09075_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_12_ ),
    .Y(_02625_)
  );
  OAI21X1 _09076_ (
    .A(_02512_),
    .B(_02620_),
    .C(_02625_),
    .Y(_02310_)
  );
  AOI22X1 _09077_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_11_ ),
    .Y(_02626_)
  );
  OAI21X1 _09078_ (
    .A(_02518_),
    .B(_02620_),
    .C(_02626_),
    .Y(_02309_)
  );
  AOI22X1 _09079_ (
    .A(_02523_),
    .B(_02619_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_10_ ),
    .Y(_02627_)
  );
  OAI21X1 _09080_ (
    .A(_02526_),
    .B(_02617_),
    .C(_02627_),
    .Y(_02308_)
  );
  AOI22X1 _09081_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_9_ ),
    .Y(_02628_)
  );
  OAI21X1 _09082_ (
    .A(_02529_),
    .B(_02620_),
    .C(_02628_),
    .Y(_02307_)
  );
  AOI22X1 _09083_ (
    .A(_02534_),
    .B(_02619_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_8_ ),
    .Y(_02629_)
  );
  OAI21X1 _09084_ (
    .A(_02537_),
    .B(_02617_),
    .C(_02629_),
    .Y(_02306_)
  );
  AOI22X1 _09085_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_7_ ),
    .Y(_02630_)
  );
  OAI21X1 _09086_ (
    .A(_02540_),
    .B(_02620_),
    .C(_02630_),
    .Y(_02305_)
  );
  AOI22X1 _09087_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_6_ ),
    .Y(_02631_)
  );
  OAI21X1 _09088_ (
    .A(_02544_),
    .B(_02620_),
    .C(_02631_),
    .Y(_02304_)
  );
  AOI22X1 _09089_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_5_ ),
    .Y(_02632_)
  );
  OAI21X1 _09090_ (
    .A(_02549_),
    .B(_02620_),
    .C(_02632_),
    .Y(_02303_)
  );
  AOI22X1 _09091_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_4_ ),
    .Y(_02633_)
  );
  OAI21X1 _09092_ (
    .A(_02553_),
    .B(_02620_),
    .C(_02633_),
    .Y(_02302_)
  );
  AOI22X1 _09093_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_3_ ),
    .Y(_02634_)
  );
  OAI21X1 _09094_ (
    .A(_02558_),
    .B(_02620_),
    .C(_02634_),
    .Y(_02301_)
  );
  AOI22X1 _09095_ (
    .A(_02562_),
    .B(_02619_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_2_ ),
    .Y(_02635_)
  );
  OAI21X1 _09096_ (
    .A(_03099_),
    .B(_02617_),
    .C(_02635_),
    .Y(_02300_)
  );
  AOI22X1 _09097_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02616_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_1_ ),
    .Y(_02636_)
  );
  OAI21X1 _09098_ (
    .A(_02566_),
    .B(_02620_),
    .C(_02636_),
    .Y(_02299_)
  );
  AOI22X1 _09099_ (
    .A(_02613_),
    .B(_02619_),
    .C(_02621_),
    .D( execution_unit_0.register_file_0.r5_0_ ),
    .Y(_02637_)
  );
  OAI21X1 _09100_ (
    .A(_03101_),
    .B(_02617_),
    .C(_02637_),
    .Y(_02298_)
  );
  AND2X1 _09101_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_6_ ),
    .Y(_02638_)
  );
  NAND2X1 _09102_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_6_ ),
    .Y(_02639_)
  );
  NAND2X1 _09103_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03124_),
    .Y(_02640_)
  );
  NOR2X1 _09104_ (
    .A(_02638_),
    .B(_02640_),
    .Y(_02641_)
  );
  OR2X1 _09105_ (
    .A(_02638_),
    .B(_02640_),
    .Y(_02642_)
  );
  AOI21X1 _09106_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03124_),
    .C(_02638_),
    .Y(_02643_)
  );
  AOI22X1 _09107_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_15_ ),
    .Y(_02644_)
  );
  OAI21X1 _09108_ (
    .A(_02491_),
    .B(_02642_),
    .C(_02644_),
    .Y(_02297_)
  );
  AOI22X1 _09109_ (
    .A(_02501_),
    .B(_02641_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_14_ ),
    .Y(_02645_)
  );
  OAI21X1 _09110_ (
    .A(_02504_),
    .B(_02639_),
    .C(_02645_),
    .Y(_02296_)
  );
  AOI22X1 _09111_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_13_ ),
    .Y(_02646_)
  );
  OAI21X1 _09112_ (
    .A(_02507_),
    .B(_02642_),
    .C(_02646_),
    .Y(_02295_)
  );
  AOI22X1 _09113_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_12_ ),
    .Y(_02647_)
  );
  OAI21X1 _09114_ (
    .A(_02512_),
    .B(_02642_),
    .C(_02647_),
    .Y(_02294_)
  );
  AOI22X1 _09115_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_11_ ),
    .Y(_02648_)
  );
  OAI21X1 _09116_ (
    .A(_02518_),
    .B(_02642_),
    .C(_02648_),
    .Y(_02293_)
  );
  AOI22X1 _09117_ (
    .A(_02523_),
    .B(_02641_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_10_ ),
    .Y(_02649_)
  );
  OAI21X1 _09118_ (
    .A(_02526_),
    .B(_02639_),
    .C(_02649_),
    .Y(_02292_)
  );
  AOI22X1 _09119_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_9_ ),
    .Y(_02650_)
  );
  OAI21X1 _09120_ (
    .A(_02529_),
    .B(_02642_),
    .C(_02650_),
    .Y(_02291_)
  );
  AOI22X1 _09121_ (
    .A(_02534_),
    .B(_02641_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_8_ ),
    .Y(_02651_)
  );
  OAI21X1 _09122_ (
    .A(_02537_),
    .B(_02639_),
    .C(_02651_),
    .Y(_02290_)
  );
  AOI22X1 _09123_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_7_ ),
    .Y(_02652_)
  );
  OAI21X1 _09124_ (
    .A(_02540_),
    .B(_02642_),
    .C(_02652_),
    .Y(_02289_)
  );
  AOI22X1 _09125_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_6_ ),
    .Y(_02653_)
  );
  OAI21X1 _09126_ (
    .A(_02544_),
    .B(_02642_),
    .C(_02653_),
    .Y(_02288_)
  );
  AOI22X1 _09127_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_5_ ),
    .Y(_02654_)
  );
  OAI21X1 _09128_ (
    .A(_02549_),
    .B(_02642_),
    .C(_02654_),
    .Y(_02287_)
  );
  AOI22X1 _09129_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_4_ ),
    .Y(_02655_)
  );
  OAI21X1 _09130_ (
    .A(_02553_),
    .B(_02642_),
    .C(_02655_),
    .Y(_02286_)
  );
  AOI22X1 _09131_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02656_)
  );
  OAI21X1 _09132_ (
    .A(_02558_),
    .B(_02642_),
    .C(_02656_),
    .Y(_02285_)
  );
  AOI22X1 _09133_ (
    .A(_02562_),
    .B(_02641_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_2_ ),
    .Y(_02657_)
  );
  OAI21X1 _09134_ (
    .A(_03099_),
    .B(_02639_),
    .C(_02657_),
    .Y(_02284_)
  );
  AOI22X1 _09135_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02638_),
    .C(_02643_),
    .D( execution_unit_0.register_file_0.r6_1_ ),
    .Y(_02658_)
  );
  OAI21X1 _09136_ (
    .A(_02566_),
    .B(_02642_),
    .C(_02658_),
    .Y(_02283_)
  );
  NAND2X1 _09137_ (
    .A( execution_unit_0.register_file_0.r6_0_ ),
    .B(_02643_),
    .Y(_02659_)
  );
  AOI22X1 _09138_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02638_),
    .C(_02641_),
    .D(_02613_),
    .Y(_02660_)
  );
  NAND2X1 _09139_ (
    .A(_02659_),
    .B(_02660_),
    .Y(_02282_)
  );
  AND2X1 _09140_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_7_ ),
    .Y(_02661_)
  );
  NAND2X1 _09141_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_7_ ),
    .Y(_02662_)
  );
  NAND2X1 _09142_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03120_),
    .Y(_02663_)
  );
  NOR2X1 _09143_ (
    .A(_02661_),
    .B(_02663_),
    .Y(_02664_)
  );
  OR2X1 _09144_ (
    .A(_02661_),
    .B(_02663_),
    .Y(_02665_)
  );
  AOI21X1 _09145_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03120_),
    .C(_02661_),
    .Y(_02666_)
  );
  AOI22X1 _09146_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_15_ ),
    .Y(_02667_)
  );
  OAI21X1 _09147_ (
    .A(_02491_),
    .B(_02665_),
    .C(_02667_),
    .Y(_02281_)
  );
  AOI22X1 _09148_ (
    .A(_02501_),
    .B(_02664_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_14_ ),
    .Y(_02668_)
  );
  OAI21X1 _09149_ (
    .A(_02504_),
    .B(_02662_),
    .C(_02668_),
    .Y(_02280_)
  );
  AOI22X1 _09150_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_13_ ),
    .Y(_02669_)
  );
  OAI21X1 _09151_ (
    .A(_02507_),
    .B(_02665_),
    .C(_02669_),
    .Y(_02279_)
  );
  AOI22X1 _09152_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_12_ ),
    .Y(_02670_)
  );
  OAI21X1 _09153_ (
    .A(_02512_),
    .B(_02665_),
    .C(_02670_),
    .Y(_02278_)
  );
  AOI22X1 _09154_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_11_ ),
    .Y(_02671_)
  );
  OAI21X1 _09155_ (
    .A(_02518_),
    .B(_02665_),
    .C(_02671_),
    .Y(_02277_)
  );
  AOI22X1 _09156_ (
    .A(_02523_),
    .B(_02664_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_10_ ),
    .Y(_02672_)
  );
  OAI21X1 _09157_ (
    .A(_02526_),
    .B(_02662_),
    .C(_02672_),
    .Y(_02276_)
  );
  AOI22X1 _09158_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_9_ ),
    .Y(_02673_)
  );
  OAI21X1 _09159_ (
    .A(_02529_),
    .B(_02665_),
    .C(_02673_),
    .Y(_02275_)
  );
  AOI22X1 _09160_ (
    .A(_02534_),
    .B(_02664_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_8_ ),
    .Y(_02674_)
  );
  OAI21X1 _09161_ (
    .A(_02537_),
    .B(_02662_),
    .C(_02674_),
    .Y(_02274_)
  );
  AOI22X1 _09162_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_7_ ),
    .Y(_02675_)
  );
  OAI21X1 _09163_ (
    .A(_02540_),
    .B(_02665_),
    .C(_02675_),
    .Y(_02273_)
  );
  AOI22X1 _09164_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_6_ ),
    .Y(_02676_)
  );
  OAI21X1 _09165_ (
    .A(_02544_),
    .B(_02665_),
    .C(_02676_),
    .Y(_02272_)
  );
  AOI22X1 _09166_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02677_)
  );
  OAI21X1 _09167_ (
    .A(_02549_),
    .B(_02665_),
    .C(_02677_),
    .Y(_02271_)
  );
  AOI22X1 _09168_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_4_ ),
    .Y(_02678_)
  );
  OAI21X1 _09169_ (
    .A(_02553_),
    .B(_02665_),
    .C(_02678_),
    .Y(_02270_)
  );
  AOI22X1 _09170_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02679_)
  );
  OAI21X1 _09171_ (
    .A(_02558_),
    .B(_02665_),
    .C(_02679_),
    .Y(_02269_)
  );
  AOI22X1 _09172_ (
    .A(_02562_),
    .B(_02664_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02680_)
  );
  OAI21X1 _09173_ (
    .A(_03099_),
    .B(_02662_),
    .C(_02680_),
    .Y(_02268_)
  );
  AOI22X1 _09174_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02661_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02681_)
  );
  OAI21X1 _09175_ (
    .A(_02566_),
    .B(_02665_),
    .C(_02681_),
    .Y(_02267_)
  );
  AOI22X1 _09176_ (
    .A(_02613_),
    .B(_02664_),
    .C(_02666_),
    .D( execution_unit_0.register_file_0.r7_0_ ),
    .Y(_02682_)
  );
  OAI21X1 _09177_ (
    .A(_03101_),
    .B(_02662_),
    .C(_02682_),
    .Y(_02266_)
  );
  AND2X1 _09178_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_8_ ),
    .Y(_02683_)
  );
  NAND2X1 _09179_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_8_ ),
    .Y(_02684_)
  );
  NAND2X1 _09180_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03116_),
    .Y(_02685_)
  );
  NOR2X1 _09181_ (
    .A(_02683_),
    .B(_02685_),
    .Y(_02686_)
  );
  OR2X1 _09182_ (
    .A(_02683_),
    .B(_02685_),
    .Y(_02687_)
  );
  AOI21X1 _09183_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03116_),
    .C(_02683_),
    .Y(_02688_)
  );
  AOI22X1 _09184_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_15_ ),
    .Y(_02689_)
  );
  OAI21X1 _09185_ (
    .A(_02491_),
    .B(_02687_),
    .C(_02689_),
    .Y(_02265_)
  );
  AOI22X1 _09186_ (
    .A(_02501_),
    .B(_02686_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_14_ ),
    .Y(_02690_)
  );
  OAI21X1 _09187_ (
    .A(_02504_),
    .B(_02684_),
    .C(_02690_),
    .Y(_02264_)
  );
  AOI22X1 _09188_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_13_ ),
    .Y(_02691_)
  );
  OAI21X1 _09189_ (
    .A(_02507_),
    .B(_02687_),
    .C(_02691_),
    .Y(_02263_)
  );
  AOI22X1 _09190_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_12_ ),
    .Y(_02692_)
  );
  OAI21X1 _09191_ (
    .A(_02512_),
    .B(_02687_),
    .C(_02692_),
    .Y(_02262_)
  );
  AOI22X1 _09192_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_11_ ),
    .Y(_02693_)
  );
  OAI21X1 _09193_ (
    .A(_02518_),
    .B(_02687_),
    .C(_02693_),
    .Y(_02261_)
  );
  AOI22X1 _09194_ (
    .A(_02523_),
    .B(_02686_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_10_ ),
    .Y(_02694_)
  );
  OAI21X1 _09195_ (
    .A(_02526_),
    .B(_02684_),
    .C(_02694_),
    .Y(_02260_)
  );
  AOI22X1 _09196_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_9_ ),
    .Y(_02695_)
  );
  OAI21X1 _09197_ (
    .A(_02529_),
    .B(_02687_),
    .C(_02695_),
    .Y(_02259_)
  );
  AOI22X1 _09198_ (
    .A(_02534_),
    .B(_02686_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_8_ ),
    .Y(_02696_)
  );
  OAI21X1 _09199_ (
    .A(_02537_),
    .B(_02684_),
    .C(_02696_),
    .Y(_02258_)
  );
  AOI22X1 _09200_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_7_ ),
    .Y(_02697_)
  );
  OAI21X1 _09201_ (
    .A(_02540_),
    .B(_02687_),
    .C(_02697_),
    .Y(_02257_)
  );
  AOI22X1 _09202_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_6_ ),
    .Y(_02698_)
  );
  OAI21X1 _09203_ (
    .A(_02544_),
    .B(_02687_),
    .C(_02698_),
    .Y(_02256_)
  );
  AOI22X1 _09204_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_5_ ),
    .Y(_02699_)
  );
  OAI21X1 _09205_ (
    .A(_02549_),
    .B(_02687_),
    .C(_02699_),
    .Y(_02255_)
  );
  AOI22X1 _09206_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_4_ ),
    .Y(_02700_)
  );
  OAI21X1 _09207_ (
    .A(_02553_),
    .B(_02687_),
    .C(_02700_),
    .Y(_02254_)
  );
  AOI22X1 _09208_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02701_)
  );
  OAI21X1 _09209_ (
    .A(_02558_),
    .B(_02687_),
    .C(_02701_),
    .Y(_02253_)
  );
  NAND2X1 _09210_ (
    .A( execution_unit_0.register_file_0.r8_2_ ),
    .B(_02688_),
    .Y(_02702_)
  );
  AOI22X1 _09211_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02683_),
    .C(_02686_),
    .D(_02562_),
    .Y(_02703_)
  );
  NAND2X1 _09212_ (
    .A(_02702_),
    .B(_02703_),
    .Y(_02252_)
  );
  AOI22X1 _09213_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02683_),
    .C(_02688_),
    .D( execution_unit_0.register_file_0.r8_1_ ),
    .Y(_02704_)
  );
  OAI21X1 _09214_ (
    .A(_02566_),
    .B(_02687_),
    .C(_02704_),
    .Y(_02251_)
  );
  NAND2X1 _09215_ (
    .A( execution_unit_0.register_file_0.r8_0_ ),
    .B(_02688_),
    .Y(_02705_)
  );
  AOI22X1 _09216_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02683_),
    .C(_02686_),
    .D(_02613_),
    .Y(_02706_)
  );
  NAND2X1 _09217_ (
    .A(_02705_),
    .B(_02706_),
    .Y(_02250_)
  );
  AND2X1 _09218_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_9_ ),
    .Y(_02707_)
  );
  NAND2X1 _09219_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_9_ ),
    .Y(_02708_)
  );
  NAND2X1 _09220_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03114_),
    .Y(_02709_)
  );
  NOR2X1 _09221_ (
    .A(_02707_),
    .B(_02709_),
    .Y(_02710_)
  );
  OR2X1 _09222_ (
    .A(_02707_),
    .B(_02709_),
    .Y(_02711_)
  );
  AOI21X1 _09223_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03114_),
    .C(_02707_),
    .Y(_02712_)
  );
  AOI22X1 _09224_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_15_ ),
    .Y(_02713_)
  );
  OAI21X1 _09225_ (
    .A(_02491_),
    .B(_02711_),
    .C(_02713_),
    .Y(_02249_)
  );
  AOI22X1 _09226_ (
    .A(_02501_),
    .B(_02710_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_14_ ),
    .Y(_02714_)
  );
  OAI21X1 _09227_ (
    .A(_02504_),
    .B(_02708_),
    .C(_02714_),
    .Y(_02248_)
  );
  AOI22X1 _09228_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_13_ ),
    .Y(_02715_)
  );
  OAI21X1 _09229_ (
    .A(_02507_),
    .B(_02711_),
    .C(_02715_),
    .Y(_02247_)
  );
  AOI22X1 _09230_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_12_ ),
    .Y(_02716_)
  );
  OAI21X1 _09231_ (
    .A(_02512_),
    .B(_02711_),
    .C(_02716_),
    .Y(_02246_)
  );
  AOI22X1 _09232_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_11_ ),
    .Y(_02717_)
  );
  OAI21X1 _09233_ (
    .A(_02518_),
    .B(_02711_),
    .C(_02717_),
    .Y(_02245_)
  );
  AOI22X1 _09234_ (
    .A(_02523_),
    .B(_02710_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_10_ ),
    .Y(_02718_)
  );
  OAI21X1 _09235_ (
    .A(_02526_),
    .B(_02708_),
    .C(_02718_),
    .Y(_02244_)
  );
  AOI22X1 _09236_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_9_ ),
    .Y(_02719_)
  );
  OAI21X1 _09237_ (
    .A(_02529_),
    .B(_02711_),
    .C(_02719_),
    .Y(_02243_)
  );
  AOI22X1 _09238_ (
    .A(_02534_),
    .B(_02710_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_8_ ),
    .Y(_02720_)
  );
  OAI21X1 _09239_ (
    .A(_02537_),
    .B(_02708_),
    .C(_02720_),
    .Y(_02242_)
  );
  AOI22X1 _09240_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_7_ ),
    .Y(_02721_)
  );
  OAI21X1 _09241_ (
    .A(_02540_),
    .B(_02711_),
    .C(_02721_),
    .Y(_02241_)
  );
  AOI22X1 _09242_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_6_ ),
    .Y(_02722_)
  );
  OAI21X1 _09243_ (
    .A(_02544_),
    .B(_02711_),
    .C(_02722_),
    .Y(_02240_)
  );
  AOI22X1 _09244_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02723_)
  );
  OAI21X1 _09245_ (
    .A(_02549_),
    .B(_02711_),
    .C(_02723_),
    .Y(_02239_)
  );
  AOI22X1 _09246_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_4_ ),
    .Y(_02724_)
  );
  OAI21X1 _09247_ (
    .A(_02553_),
    .B(_02711_),
    .C(_02724_),
    .Y(_02238_)
  );
  AOI22X1 _09248_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_3_ ),
    .Y(_02725_)
  );
  OAI21X1 _09249_ (
    .A(_02558_),
    .B(_02711_),
    .C(_02725_),
    .Y(_02237_)
  );
  AOI22X1 _09250_ (
    .A(_02562_),
    .B(_02710_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_2_ ),
    .Y(_02726_)
  );
  OAI21X1 _09251_ (
    .A(_03099_),
    .B(_02708_),
    .C(_02726_),
    .Y(_02236_)
  );
  AOI22X1 _09252_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02707_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_1_ ),
    .Y(_02727_)
  );
  OAI21X1 _09253_ (
    .A(_02566_),
    .B(_02711_),
    .C(_02727_),
    .Y(_02235_)
  );
  AOI22X1 _09254_ (
    .A(_02613_),
    .B(_02710_),
    .C(_02712_),
    .D( execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02728_)
  );
  OAI21X1 _09255_ (
    .A(_03101_),
    .B(_02708_),
    .C(_02728_),
    .Y(_02234_)
  );
  AND2X1 _09256_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_10_ ),
    .Y(_02729_)
  );
  NAND2X1 _09257_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_10_ ),
    .Y(_02730_)
  );
  NAND2X1 _09258_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03115_),
    .Y(_02731_)
  );
  NOR2X1 _09259_ (
    .A(_02729_),
    .B(_02731_),
    .Y(_02732_)
  );
  OR2X1 _09260_ (
    .A(_02729_),
    .B(_02731_),
    .Y(_02733_)
  );
  AOI21X1 _09261_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03115_),
    .C(_02729_),
    .Y(_02734_)
  );
  AOI22X1 _09262_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02735_)
  );
  OAI21X1 _09263_ (
    .A(_02491_),
    .B(_02733_),
    .C(_02735_),
    .Y(_02233_)
  );
  AOI22X1 _09264_ (
    .A(_02501_),
    .B(_02732_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_14_ ),
    .Y(_02736_)
  );
  OAI21X1 _09265_ (
    .A(_02504_),
    .B(_02730_),
    .C(_02736_),
    .Y(_02232_)
  );
  AOI22X1 _09266_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_13_ ),
    .Y(_02737_)
  );
  OAI21X1 _09267_ (
    .A(_02507_),
    .B(_02733_),
    .C(_02737_),
    .Y(_02231_)
  );
  AOI22X1 _09268_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_12_ ),
    .Y(_02738_)
  );
  OAI21X1 _09269_ (
    .A(_02512_),
    .B(_02733_),
    .C(_02738_),
    .Y(_02230_)
  );
  AOI22X1 _09270_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_11_ ),
    .Y(_02739_)
  );
  OAI21X1 _09271_ (
    .A(_02518_),
    .B(_02733_),
    .C(_02739_),
    .Y(_02229_)
  );
  AOI22X1 _09272_ (
    .A(_02523_),
    .B(_02732_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_10_ ),
    .Y(_02740_)
  );
  OAI21X1 _09273_ (
    .A(_02526_),
    .B(_02730_),
    .C(_02740_),
    .Y(_02228_)
  );
  AOI22X1 _09274_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_9_ ),
    .Y(_02741_)
  );
  OAI21X1 _09275_ (
    .A(_02529_),
    .B(_02733_),
    .C(_02741_),
    .Y(_02227_)
  );
  AOI22X1 _09276_ (
    .A(_02534_),
    .B(_02732_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_8_ ),
    .Y(_02742_)
  );
  OAI21X1 _09277_ (
    .A(_02537_),
    .B(_02730_),
    .C(_02742_),
    .Y(_02226_)
  );
  AOI22X1 _09278_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_7_ ),
    .Y(_02743_)
  );
  OAI21X1 _09279_ (
    .A(_02540_),
    .B(_02733_),
    .C(_02743_),
    .Y(_02225_)
  );
  AOI22X1 _09280_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_6_ ),
    .Y(_02744_)
  );
  OAI21X1 _09281_ (
    .A(_02544_),
    .B(_02733_),
    .C(_02744_),
    .Y(_02224_)
  );
  AOI22X1 _09282_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_5_ ),
    .Y(_02745_)
  );
  OAI21X1 _09283_ (
    .A(_02549_),
    .B(_02733_),
    .C(_02745_),
    .Y(_02223_)
  );
  AOI22X1 _09284_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_4_ ),
    .Y(_02746_)
  );
  OAI21X1 _09285_ (
    .A(_02553_),
    .B(_02733_),
    .C(_02746_),
    .Y(_02222_)
  );
  AOI22X1 _09286_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_3_ ),
    .Y(_02747_)
  );
  OAI21X1 _09287_ (
    .A(_02558_),
    .B(_02733_),
    .C(_02747_),
    .Y(_02221_)
  );
  NAND2X1 _09288_ (
    .A( execution_unit_0.register_file_0.r10_2_ ),
    .B(_02734_),
    .Y(_02748_)
  );
  AOI22X1 _09289_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02729_),
    .C(_02732_),
    .D(_02562_),
    .Y(_02749_)
  );
  NAND2X1 _09290_ (
    .A(_02748_),
    .B(_02749_),
    .Y(_02220_)
  );
  AOI22X1 _09291_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02729_),
    .C(_02734_),
    .D( execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02750_)
  );
  OAI21X1 _09292_ (
    .A(_02566_),
    .B(_02733_),
    .C(_02750_),
    .Y(_02219_)
  );
  NAND2X1 _09293_ (
    .A( execution_unit_0.register_file_0.r10_0_ ),
    .B(_02734_),
    .Y(_02751_)
  );
  AOI22X1 _09294_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02729_),
    .C(_02732_),
    .D(_02613_),
    .Y(_02752_)
  );
  NAND2X1 _09295_ (
    .A(_02751_),
    .B(_02752_),
    .Y(_02218_)
  );
  AND2X1 _09296_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_11_ ),
    .Y(_02753_)
  );
  NAND2X1 _09297_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_11_ ),
    .Y(_02754_)
  );
  NAND2X1 _09298_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03112_),
    .Y(_02755_)
  );
  NOR2X1 _09299_ (
    .A(_02753_),
    .B(_02755_),
    .Y(_02756_)
  );
  OR2X1 _09300_ (
    .A(_02753_),
    .B(_02755_),
    .Y(_02757_)
  );
  AOI21X1 _09301_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03112_),
    .C(_02753_),
    .Y(_02758_)
  );
  AOI22X1 _09302_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_15_ ),
    .Y(_02759_)
  );
  OAI21X1 _09303_ (
    .A(_02491_),
    .B(_02757_),
    .C(_02759_),
    .Y(_02217_)
  );
  AOI22X1 _09304_ (
    .A(_02501_),
    .B(_02756_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_14_ ),
    .Y(_02760_)
  );
  OAI21X1 _09305_ (
    .A(_02504_),
    .B(_02754_),
    .C(_02760_),
    .Y(_02216_)
  );
  AOI22X1 _09306_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_13_ ),
    .Y(_02761_)
  );
  OAI21X1 _09307_ (
    .A(_02507_),
    .B(_02757_),
    .C(_02761_),
    .Y(_02215_)
  );
  AOI22X1 _09308_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_12_ ),
    .Y(_02762_)
  );
  OAI21X1 _09309_ (
    .A(_02512_),
    .B(_02757_),
    .C(_02762_),
    .Y(_02214_)
  );
  AOI22X1 _09310_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_11_ ),
    .Y(_02763_)
  );
  OAI21X1 _09311_ (
    .A(_02518_),
    .B(_02757_),
    .C(_02763_),
    .Y(_02213_)
  );
  AOI22X1 _09312_ (
    .A(_02523_),
    .B(_02756_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_10_ ),
    .Y(_02764_)
  );
  OAI21X1 _09313_ (
    .A(_02526_),
    .B(_02754_),
    .C(_02764_),
    .Y(_02212_)
  );
  AOI22X1 _09314_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_9_ ),
    .Y(_02765_)
  );
  OAI21X1 _09315_ (
    .A(_02529_),
    .B(_02757_),
    .C(_02765_),
    .Y(_02211_)
  );
  AOI22X1 _09316_ (
    .A(_02534_),
    .B(_02756_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_8_ ),
    .Y(_02766_)
  );
  OAI21X1 _09317_ (
    .A(_02537_),
    .B(_02754_),
    .C(_02766_),
    .Y(_02210_)
  );
  AOI22X1 _09318_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_7_ ),
    .Y(_02767_)
  );
  OAI21X1 _09319_ (
    .A(_02540_),
    .B(_02757_),
    .C(_02767_),
    .Y(_02209_)
  );
  AOI22X1 _09320_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_6_ ),
    .Y(_02768_)
  );
  OAI21X1 _09321_ (
    .A(_02544_),
    .B(_02757_),
    .C(_02768_),
    .Y(_02208_)
  );
  AOI22X1 _09322_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_5_ ),
    .Y(_02769_)
  );
  OAI21X1 _09323_ (
    .A(_02549_),
    .B(_02757_),
    .C(_02769_),
    .Y(_02207_)
  );
  AOI22X1 _09324_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02770_)
  );
  OAI21X1 _09325_ (
    .A(_02553_),
    .B(_02757_),
    .C(_02770_),
    .Y(_02206_)
  );
  AOI22X1 _09326_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_3_ ),
    .Y(_02771_)
  );
  OAI21X1 _09327_ (
    .A(_02558_),
    .B(_02757_),
    .C(_02771_),
    .Y(_02205_)
  );
  AOI22X1 _09328_ (
    .A(_02562_),
    .B(_02756_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_2_ ),
    .Y(_02772_)
  );
  OAI21X1 _09329_ (
    .A(_03099_),
    .B(_02754_),
    .C(_02772_),
    .Y(_02204_)
  );
  AOI22X1 _09330_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02753_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02773_)
  );
  OAI21X1 _09331_ (
    .A(_02566_),
    .B(_02757_),
    .C(_02773_),
    .Y(_02203_)
  );
  AOI22X1 _09332_ (
    .A(_02613_),
    .B(_02756_),
    .C(_02758_),
    .D( execution_unit_0.register_file_0.r11_0_ ),
    .Y(_02774_)
  );
  OAI21X1 _09333_ (
    .A(_03101_),
    .B(_02754_),
    .C(_02774_),
    .Y(_02202_)
  );
  AND2X1 _09334_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_02775_)
  );
  NAND2X1 _09335_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_02776_)
  );
  NAND2X1 _09336_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03125_),
    .Y(_02777_)
  );
  NOR2X1 _09337_ (
    .A(_02775_),
    .B(_02777_),
    .Y(_02778_)
  );
  OR2X1 _09338_ (
    .A(_02775_),
    .B(_02777_),
    .Y(_02779_)
  );
  AOI21X1 _09339_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03125_),
    .C(_02775_),
    .Y(_02780_)
  );
  AOI22X1 _09340_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_15_ ),
    .Y(_02781_)
  );
  OAI21X1 _09341_ (
    .A(_02491_),
    .B(_02779_),
    .C(_02781_),
    .Y(_02201_)
  );
  AOI22X1 _09342_ (
    .A(_02501_),
    .B(_02778_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_02782_)
  );
  OAI21X1 _09343_ (
    .A(_02504_),
    .B(_02776_),
    .C(_02782_),
    .Y(_02200_)
  );
  AOI22X1 _09344_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_13_ ),
    .Y(_02783_)
  );
  OAI21X1 _09345_ (
    .A(_02507_),
    .B(_02779_),
    .C(_02783_),
    .Y(_02199_)
  );
  AOI22X1 _09346_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_12_ ),
    .Y(_02784_)
  );
  OAI21X1 _09347_ (
    .A(_02512_),
    .B(_02779_),
    .C(_02784_),
    .Y(_02198_)
  );
  AOI22X1 _09348_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_11_ ),
    .Y(_02785_)
  );
  OAI21X1 _09349_ (
    .A(_02518_),
    .B(_02779_),
    .C(_02785_),
    .Y(_02197_)
  );
  AOI22X1 _09350_ (
    .A(_02523_),
    .B(_02778_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_10_ ),
    .Y(_02786_)
  );
  OAI21X1 _09351_ (
    .A(_02526_),
    .B(_02776_),
    .C(_02786_),
    .Y(_02196_)
  );
  AOI22X1 _09352_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_9_ ),
    .Y(_02787_)
  );
  OAI21X1 _09353_ (
    .A(_02529_),
    .B(_02779_),
    .C(_02787_),
    .Y(_02195_)
  );
  AOI22X1 _09354_ (
    .A(_02534_),
    .B(_02778_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_8_ ),
    .Y(_02788_)
  );
  OAI21X1 _09355_ (
    .A(_02537_),
    .B(_02776_),
    .C(_02788_),
    .Y(_02194_)
  );
  AOI22X1 _09356_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_7_ ),
    .Y(_02789_)
  );
  OAI21X1 _09357_ (
    .A(_02540_),
    .B(_02779_),
    .C(_02789_),
    .Y(_02193_)
  );
  AOI22X1 _09358_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_6_ ),
    .Y(_02790_)
  );
  OAI21X1 _09359_ (
    .A(_02544_),
    .B(_02779_),
    .C(_02790_),
    .Y(_02192_)
  );
  AOI22X1 _09360_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02791_)
  );
  OAI21X1 _09361_ (
    .A(_02549_),
    .B(_02779_),
    .C(_02791_),
    .Y(_02191_)
  );
  AOI22X1 _09362_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02792_)
  );
  OAI21X1 _09363_ (
    .A(_02553_),
    .B(_02779_),
    .C(_02792_),
    .Y(_02190_)
  );
  AOI22X1 _09364_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_3_ ),
    .Y(_02793_)
  );
  OAI21X1 _09365_ (
    .A(_02558_),
    .B(_02779_),
    .C(_02793_),
    .Y(_02189_)
  );
  NAND2X1 _09366_ (
    .A( execution_unit_0.register_file_0.r12_2_ ),
    .B(_02780_),
    .Y(_02794_)
  );
  AOI22X1 _09367_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02775_),
    .C(_02778_),
    .D(_02562_),
    .Y(_02795_)
  );
  NAND2X1 _09368_ (
    .A(_02794_),
    .B(_02795_),
    .Y(_02188_)
  );
  AOI22X1 _09369_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02775_),
    .C(_02780_),
    .D( execution_unit_0.register_file_0.r12_1_ ),
    .Y(_02796_)
  );
  OAI21X1 _09370_ (
    .A(_02566_),
    .B(_02779_),
    .C(_02796_),
    .Y(_02187_)
  );
  NAND2X1 _09371_ (
    .A( execution_unit_0.register_file_0.r12_0_ ),
    .B(_02780_),
    .Y(_02797_)
  );
  AOI22X1 _09372_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02775_),
    .C(_02778_),
    .D(_02613_),
    .Y(_02798_)
  );
  NAND2X1 _09373_ (
    .A(_02797_),
    .B(_02798_),
    .Y(_02186_)
  );
  AND2X1 _09374_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_02799_)
  );
  NAND2X1 _09375_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_02800_)
  );
  NAND2X1 _09376_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03111_),
    .Y(_02801_)
  );
  NOR2X1 _09377_ (
    .A(_02799_),
    .B(_02801_),
    .Y(_02802_)
  );
  OR2X1 _09378_ (
    .A(_02799_),
    .B(_02801_),
    .Y(_02803_)
  );
  AOI21X1 _09379_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03111_),
    .C(_02799_),
    .Y(_02804_)
  );
  AOI22X1 _09380_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_15_ ),
    .Y(_02805_)
  );
  OAI21X1 _09381_ (
    .A(_02491_),
    .B(_02803_),
    .C(_02805_),
    .Y(_02185_)
  );
  AOI22X1 _09382_ (
    .A(_02501_),
    .B(_02802_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_14_ ),
    .Y(_02806_)
  );
  OAI21X1 _09383_ (
    .A(_02504_),
    .B(_02800_),
    .C(_02806_),
    .Y(_02184_)
  );
  AOI22X1 _09384_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_13_ ),
    .Y(_02807_)
  );
  OAI21X1 _09385_ (
    .A(_02507_),
    .B(_02803_),
    .C(_02807_),
    .Y(_02183_)
  );
  AOI22X1 _09386_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_12_ ),
    .Y(_02808_)
  );
  OAI21X1 _09387_ (
    .A(_02512_),
    .B(_02803_),
    .C(_02808_),
    .Y(_02182_)
  );
  AOI22X1 _09388_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_11_ ),
    .Y(_02809_)
  );
  OAI21X1 _09389_ (
    .A(_02518_),
    .B(_02803_),
    .C(_02809_),
    .Y(_02181_)
  );
  AOI22X1 _09390_ (
    .A(_02523_),
    .B(_02802_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_10_ ),
    .Y(_02810_)
  );
  OAI21X1 _09391_ (
    .A(_02526_),
    .B(_02800_),
    .C(_02810_),
    .Y(_02180_)
  );
  AOI22X1 _09392_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_9_ ),
    .Y(_02811_)
  );
  OAI21X1 _09393_ (
    .A(_02529_),
    .B(_02803_),
    .C(_02811_),
    .Y(_02179_)
  );
  AOI22X1 _09394_ (
    .A(_02534_),
    .B(_02802_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_8_ ),
    .Y(_02812_)
  );
  OAI21X1 _09395_ (
    .A(_02537_),
    .B(_02800_),
    .C(_02812_),
    .Y(_02178_)
  );
  AOI22X1 _09396_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_7_ ),
    .Y(_02813_)
  );
  OAI21X1 _09397_ (
    .A(_02540_),
    .B(_02803_),
    .C(_02813_),
    .Y(_02177_)
  );
  AOI22X1 _09398_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_6_ ),
    .Y(_02814_)
  );
  OAI21X1 _09399_ (
    .A(_02544_),
    .B(_02803_),
    .C(_02814_),
    .Y(_02176_)
  );
  AOI22X1 _09400_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_5_ ),
    .Y(_02815_)
  );
  OAI21X1 _09401_ (
    .A(_02549_),
    .B(_02803_),
    .C(_02815_),
    .Y(_02175_)
  );
  AOI22X1 _09402_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_4_ ),
    .Y(_02816_)
  );
  OAI21X1 _09403_ (
    .A(_02553_),
    .B(_02803_),
    .C(_02816_),
    .Y(_02174_)
  );
  AOI22X1 _09404_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_3_ ),
    .Y(_02817_)
  );
  OAI21X1 _09405_ (
    .A(_02558_),
    .B(_02803_),
    .C(_02817_),
    .Y(_02173_)
  );
  NAND2X1 _09406_ (
    .A( execution_unit_0.register_file_0.r13_2_ ),
    .B(_02804_),
    .Y(_02818_)
  );
  AOI22X1 _09407_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02799_),
    .C(_02802_),
    .D(_02562_),
    .Y(_02819_)
  );
  NAND2X1 _09408_ (
    .A(_02818_),
    .B(_02819_),
    .Y(_02172_)
  );
  AOI22X1 _09409_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02799_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_1_ ),
    .Y(_02820_)
  );
  OAI21X1 _09410_ (
    .A(_02566_),
    .B(_02803_),
    .C(_02820_),
    .Y(_02171_)
  );
  AOI22X1 _09411_ (
    .A(_02613_),
    .B(_02802_),
    .C(_02804_),
    .D( execution_unit_0.register_file_0.r13_0_ ),
    .Y(_02821_)
  );
  OAI21X1 _09412_ (
    .A(_03101_),
    .B(_02800_),
    .C(_02821_),
    .Y(_02170_)
  );
  AND2X1 _09413_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_14_ ),
    .Y(_02822_)
  );
  NAND2X1 _09414_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_14_ ),
    .Y(_02823_)
  );
  NAND2X1 _09415_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03123_),
    .Y(_02824_)
  );
  NOR2X1 _09416_ (
    .A(_02822_),
    .B(_02824_),
    .Y(_02825_)
  );
  OR2X1 _09417_ (
    .A(_02822_),
    .B(_02824_),
    .Y(_02826_)
  );
  AOI21X1 _09418_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03123_),
    .C(_02822_),
    .Y(_02827_)
  );
  AOI22X1 _09419_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_15_ ),
    .Y(_02828_)
  );
  OAI21X1 _09420_ (
    .A(_02491_),
    .B(_02826_),
    .C(_02828_),
    .Y(_02169_)
  );
  AOI22X1 _09421_ (
    .A(_02501_),
    .B(_02825_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_14_ ),
    .Y(_02829_)
  );
  OAI21X1 _09422_ (
    .A(_02504_),
    .B(_02823_),
    .C(_02829_),
    .Y(_02168_)
  );
  AOI22X1 _09423_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_13_ ),
    .Y(_02830_)
  );
  OAI21X1 _09424_ (
    .A(_02507_),
    .B(_02826_),
    .C(_02830_),
    .Y(_02167_)
  );
  AOI22X1 _09425_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_12_ ),
    .Y(_02831_)
  );
  OAI21X1 _09426_ (
    .A(_02512_),
    .B(_02826_),
    .C(_02831_),
    .Y(_02166_)
  );
  AOI22X1 _09427_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_11_ ),
    .Y(_02832_)
  );
  OAI21X1 _09428_ (
    .A(_02518_),
    .B(_02826_),
    .C(_02832_),
    .Y(_02165_)
  );
  AOI22X1 _09429_ (
    .A(_02523_),
    .B(_02825_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_10_ ),
    .Y(_02833_)
  );
  OAI21X1 _09430_ (
    .A(_02526_),
    .B(_02823_),
    .C(_02833_),
    .Y(_02164_)
  );
  AOI22X1 _09431_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_9_ ),
    .Y(_02834_)
  );
  OAI21X1 _09432_ (
    .A(_02529_),
    .B(_02826_),
    .C(_02834_),
    .Y(_02163_)
  );
  AOI22X1 _09433_ (
    .A(_02534_),
    .B(_02825_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_8_ ),
    .Y(_02835_)
  );
  OAI21X1 _09434_ (
    .A(_02537_),
    .B(_02823_),
    .C(_02835_),
    .Y(_02162_)
  );
  AOI22X1 _09435_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_7_ ),
    .Y(_02836_)
  );
  OAI21X1 _09436_ (
    .A(_02540_),
    .B(_02826_),
    .C(_02836_),
    .Y(_02161_)
  );
  AOI22X1 _09437_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_6_ ),
    .Y(_02837_)
  );
  OAI21X1 _09438_ (
    .A(_02544_),
    .B(_02826_),
    .C(_02837_),
    .Y(_02160_)
  );
  AOI22X1 _09439_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_5_ ),
    .Y(_02838_)
  );
  OAI21X1 _09440_ (
    .A(_02549_),
    .B(_02826_),
    .C(_02838_),
    .Y(_02159_)
  );
  AOI22X1 _09441_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_4_ ),
    .Y(_02839_)
  );
  OAI21X1 _09442_ (
    .A(_02553_),
    .B(_02826_),
    .C(_02839_),
    .Y(_02158_)
  );
  AOI22X1 _09443_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_3_ ),
    .Y(_02840_)
  );
  OAI21X1 _09444_ (
    .A(_02558_),
    .B(_02826_),
    .C(_02840_),
    .Y(_02157_)
  );
  AOI22X1 _09445_ (
    .A(_02562_),
    .B(_02825_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_2_ ),
    .Y(_02841_)
  );
  OAI21X1 _09446_ (
    .A(_03099_),
    .B(_02823_),
    .C(_02841_),
    .Y(_02156_)
  );
  AOI22X1 _09447_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02822_),
    .C(_02827_),
    .D( execution_unit_0.register_file_0.r14_1_ ),
    .Y(_02842_)
  );
  OAI21X1 _09448_ (
    .A(_02566_),
    .B(_02826_),
    .C(_02842_),
    .Y(_02155_)
  );
  NAND2X1 _09449_ (
    .A( execution_unit_0.register_file_0.r14_0_ ),
    .B(_02827_),
    .Y(_02843_)
  );
  AOI22X1 _09450_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02822_),
    .C(_02825_),
    .D(_02613_),
    .Y(_02844_)
  );
  NAND2X1 _09451_ (
    .A(_02843_),
    .B(_02844_),
    .Y(_02154_)
  );
  AND2X1 _09452_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_15_ ),
    .Y(_02845_)
  );
  NAND2X1 _09453_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_15_ ),
    .Y(_02846_)
  );
  NAND2X1 _09454_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03119_),
    .Y(_02847_)
  );
  NOR2X1 _09455_ (
    .A(_02845_),
    .B(_02847_),
    .Y(_02848_)
  );
  OR2X1 _09456_ (
    .A(_02845_),
    .B(_02847_),
    .Y(_02849_)
  );
  AOI21X1 _09457_ (
    .A( execution_unit_0.reg_incr ),
    .B(_03119_),
    .C(_02845_),
    .Y(_02850_)
  );
  AOI22X1 _09458_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_15_ ),
    .Y(_02851_)
  );
  OAI21X1 _09459_ (
    .A(_02491_),
    .B(_02849_),
    .C(_02851_),
    .Y(_02153_)
  );
  AOI22X1 _09460_ (
    .A(_02501_),
    .B(_02848_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_14_ ),
    .Y(_02852_)
  );
  OAI21X1 _09461_ (
    .A(_02504_),
    .B(_02846_),
    .C(_02852_),
    .Y(_02152_)
  );
  AOI22X1 _09462_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_13_ ),
    .Y(_02853_)
  );
  OAI21X1 _09463_ (
    .A(_02507_),
    .B(_02849_),
    .C(_02853_),
    .Y(_02151_)
  );
  AOI22X1 _09464_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_12_ ),
    .Y(_02854_)
  );
  OAI21X1 _09465_ (
    .A(_02512_),
    .B(_02849_),
    .C(_02854_),
    .Y(_02150_)
  );
  AOI22X1 _09466_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_11_ ),
    .Y(_02855_)
  );
  OAI21X1 _09467_ (
    .A(_02518_),
    .B(_02849_),
    .C(_02855_),
    .Y(_02149_)
  );
  AOI22X1 _09468_ (
    .A(_02523_),
    .B(_02848_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_10_ ),
    .Y(_02856_)
  );
  OAI21X1 _09469_ (
    .A(_02526_),
    .B(_02846_),
    .C(_02856_),
    .Y(_02148_)
  );
  AOI22X1 _09470_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_9_ ),
    .Y(_02857_)
  );
  OAI21X1 _09471_ (
    .A(_02529_),
    .B(_02849_),
    .C(_02857_),
    .Y(_02147_)
  );
  AOI22X1 _09472_ (
    .A(_02534_),
    .B(_02848_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_8_ ),
    .Y(_02858_)
  );
  OAI21X1 _09473_ (
    .A(_02537_),
    .B(_02846_),
    .C(_02858_),
    .Y(_02146_)
  );
  AOI22X1 _09474_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_7_ ),
    .Y(_02859_)
  );
  OAI21X1 _09475_ (
    .A(_02540_),
    .B(_02849_),
    .C(_02859_),
    .Y(_02145_)
  );
  AOI22X1 _09476_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_6_ ),
    .Y(_02860_)
  );
  OAI21X1 _09477_ (
    .A(_02544_),
    .B(_02849_),
    .C(_02860_),
    .Y(_02144_)
  );
  AOI22X1 _09478_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_5_ ),
    .Y(_02861_)
  );
  OAI21X1 _09479_ (
    .A(_02549_),
    .B(_02849_),
    .C(_02861_),
    .Y(_02143_)
  );
  AOI22X1 _09480_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_4_ ),
    .Y(_02862_)
  );
  OAI21X1 _09481_ (
    .A(_02553_),
    .B(_02849_),
    .C(_02862_),
    .Y(_02142_)
  );
  AOI22X1 _09482_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_3_ ),
    .Y(_02863_)
  );
  OAI21X1 _09483_ (
    .A(_02558_),
    .B(_02849_),
    .C(_02863_),
    .Y(_02141_)
  );
  AOI22X1 _09484_ (
    .A(_02562_),
    .B(_02848_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_2_ ),
    .Y(_02864_)
  );
  OAI21X1 _09485_ (
    .A(_03099_),
    .B(_02846_),
    .C(_02864_),
    .Y(_02140_)
  );
  AOI22X1 _09486_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02845_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_1_ ),
    .Y(_02865_)
  );
  OAI21X1 _09487_ (
    .A(_02566_),
    .B(_02849_),
    .C(_02865_),
    .Y(_02139_)
  );
  AOI22X1 _09488_ (
    .A(_02613_),
    .B(_02848_),
    .C(_02850_),
    .D( execution_unit_0.register_file_0.r15_0_ ),
    .Y(_02866_)
  );
  OAI21X1 _09489_ (
    .A(_03101_),
    .B(_02846_),
    .C(_02866_),
    .Y(_02138_)
  );
  NAND2X1 _09490_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B(_02570_),
    .Y(_02867_)
  );
  OAI21X1 _09491_ (
    .A(_02537_),
    .B(_02570_),
    .C(_02867_),
    .Y(_02868_)
  );
  OAI21X1 _09492_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_02868_),
    .C(_03105_),
    .Y(_02869_)
  );
  AOI21X1 _09493_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_03110_),
    .C(_02869_),
    .Y(_02137_)
  );
  AND2X1 _09494_ (
    .A(_03105_),
    .B(_02570_),
    .Y(_02870_)
  );
  NAND2X1 _09495_ (
    .A( clock_module_0.scg1 ),
    .B(_02870_),
    .Y(_02871_)
  );
  NAND2X1 _09496_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_03105_),
    .Y(_02872_)
  );
  OAI21X1 _09497_ (
    .A(_02570_),
    .B(_02872_),
    .C(_02871_),
    .Y(_02136_)
  );
  NAND2X1 _09498_ (
    .A( clock_module_0.oscoff ),
    .B(_02870_),
    .Y(_02873_)
  );
  NAND2X1 _09499_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_03105_),
    .Y(_02874_)
  );
  OAI21X1 _09500_ (
    .A(_02570_),
    .B(_02874_),
    .C(_02873_),
    .Y(_02135_)
  );
  NAND2X1 _09501_ (
    .A( execution_unit_0.gie ),
    .B(_02870_),
    .Y(_02875_)
  );
  NAND2X1 _09502_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_03105_),
    .Y(_02876_)
  );
  OAI21X1 _09503_ (
    .A(_02570_),
    .B(_02876_),
    .C(_02875_),
    .Y(_02134_)
  );
  NOR2X1 _09504_ (
    .A(_03099_),
    .B(_02570_),
    .Y(_02877_)
  );
  AOI22X1 _09505_ (
    .A( execution_unit_0.alu_0.status_2_ ),
    .B(_02870_),
    .C(_02877_),
    .D(_03105_),
    .Y(_02878_)
  );
  NAND3X1 _09506_ (
    .A(_03105_),
    .B( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .C( execution_unit_0.alu_0.N ),
    .Y(_02879_)
  );
  OAI21X1 _09507_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_02878_),
    .C(_02879_),
    .Y(_02133_)
  );
  NOR2X1 _09508_ (
    .A(_03100_),
    .B(_02570_),
    .Y(_02880_)
  );
  AOI22X1 _09509_ (
    .A( execution_unit_0.alu_0.status_1_ ),
    .B(_02870_),
    .C(_02880_),
    .D(_03105_),
    .Y(_02881_)
  );
  NAND3X1 _09510_ (
    .A(_03105_),
    .B( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .C( execution_unit_0.alu_0.Z ),
    .Y(_02882_)
  );
  OAI21X1 _09511_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_02881_),
    .C(_02882_),
    .Y(_02132_)
  );
  OAI21X1 _09512_ (
    .A(_03097_),
    .B(_02570_),
    .C(_03109_),
    .Y( clock_module_0.UNUSED_cpuoff )
  );
  MUX2X1 _09513_ (
    .A( execution_unit_0.register_file_0.r2_4_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .S(_02570_),
    .Y(_02883_)
  );
  NOR2X1 _09514_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_02883_),
    .Y(_01900_)
  );
  AOI21X1 _09515_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_0_ ),
    .C( execution_unit_0.reg_pc_call ),
    .Y(_02884_)
  );
  INVX1 _09516_ (
    .A(_02884_),
    .Y( execution_unit_0.pc_sw_wr )
  );
  NAND2X1 _09517_ (
    .A( execution_unit_0.register_file_0.r13_0_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_02885_)
  );
  AOI22X1 _09518_ (
    .A( execution_unit_0.register_file_0.r12_0_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_0_ ),
    .Y(_02886_)
  );
  AOI22X1 _09519_ (
    .A( execution_unit_0.register_file_0.r6_0_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_0_ ),
    .Y(_02887_)
  );
  AOI22X1 _09520_ (
    .A( execution_unit_0.register_file_0.r7_0_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_0_ ),
    .Y(_02888_)
  );
  NAND2X1 _09521_ (
    .A(_02885_),
    .B(_02888_),
    .Y(_02889_)
  );
  AOI21X1 _09522_ (
    .A( execution_unit_0.register_file_0.r10_0_ ),
    .B( execution_unit_0.inst_dest_10_ ),
    .C(_02889_),
    .Y(_02890_)
  );
  AND2X1 _09523_ (
    .A(_02886_),
    .B(_02887_),
    .Y(_02891_)
  );
  AOI22X1 _09524_ (
    .A( execution_unit_0.register_file_0.r9_0_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_0_ ),
    .Y(_02892_)
  );
  AOI22X1 _09525_ (
    .A( execution_unit_0.register_file_0.r15_0_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( dbg_0.UNUSED_pc_0_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02893_)
  );
  AOI22X1 _09526_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_0_ ),
    .Y(_02894_)
  );
  NAND3X1 _09527_ (
    .A(_02892_),
    .B(_02893_),
    .C(_02894_),
    .Y(_02895_)
  );
  AOI21X1 _09528_ (
    .A( execution_unit_0.register_file_0.r8_0_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C(_02895_),
    .Y(_02896_)
  );
  NAND3X1 _09529_ (
    .A(_02890_),
    .B(_02891_),
    .C(_02896_),
    .Y( dbg_0.dbg_reg_din_0_ )
  );
  AOI22X1 _09530_ (
    .A( execution_unit_0.register_file_0.r6_1_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02897_)
  );
  AOI22X1 _09531_ (
    .A( execution_unit_0.alu_0.status_1_ ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( dbg_0.UNUSED_pc_1_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02898_)
  );
  NAND2X1 _09532_ (
    .A(_02897_),
    .B(_02898_),
    .Y(_02899_)
  );
  AOI22X1 _09533_ (
    .A( execution_unit_0.register_file_0.r13_1_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_1_ ),
    .Y(_02900_)
  );
  AOI22X1 _09534_ (
    .A( execution_unit_0.register_file_0.r4_1_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02901_)
  );
  NAND2X1 _09535_ (
    .A(_02900_),
    .B(_02901_),
    .Y(_02902_)
  );
  NOR2X1 _09536_ (
    .A(_02899_),
    .B(_02902_),
    .Y(_02903_)
  );
  AOI22X1 _09537_ (
    .A( execution_unit_0.register_file_0.r1_1_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_1_ ),
    .Y(_02904_)
  );
  AOI22X1 _09538_ (
    .A( execution_unit_0.register_file_0.r8_1_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_15_ ),
    .D( execution_unit_0.register_file_0.r15_1_ ),
    .Y(_02905_)
  );
  NAND2X1 _09539_ (
    .A(_02904_),
    .B(_02905_),
    .Y(_02906_)
  );
  AOI22X1 _09540_ (
    .A( execution_unit_0.register_file_0.r9_1_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_1_ ),
    .Y(_02907_)
  );
  AOI22X1 _09541_ (
    .A( execution_unit_0.register_file_0.r7_1_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_1_ ),
    .Y(_02908_)
  );
  NAND2X1 _09542_ (
    .A(_02907_),
    .B(_02908_),
    .Y(_02909_)
  );
  NOR2X1 _09543_ (
    .A(_02906_),
    .B(_02909_),
    .Y(_02910_)
  );
  NAND2X1 _09544_ (
    .A(_02903_),
    .B(_02910_),
    .Y( dbg_0.dbg_reg_din_1_ )
  );
  AOI22X1 _09545_ (
    .A( execution_unit_0.register_file_0.r12_2_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_2_ ),
    .Y(_02911_)
  );
  AOI22X1 _09546_ (
    .A( execution_unit_0.register_file_0.r11_2_ ),
    .B( execution_unit_0.inst_dest_11_ ),
    .C( dbg_0.UNUSED_pc_2_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02912_)
  );
  NAND2X1 _09547_ (
    .A(_02911_),
    .B(_02912_),
    .Y(_02913_)
  );
  AOI22X1 _09548_ (
    .A( execution_unit_0.register_file_0.r1_2_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_2_ ),
    .Y(_02914_)
  );
  AOI22X1 _09549_ (
    .A( execution_unit_0.register_file_0.r8_2_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_7_ ),
    .D( execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02915_)
  );
  NAND2X1 _09550_ (
    .A(_02914_),
    .B(_02915_),
    .Y(_02916_)
  );
  NOR2X1 _09551_ (
    .A(_02913_),
    .B(_02916_),
    .Y(_02917_)
  );
  AOI22X1 _09552_ (
    .A( execution_unit_0.register_file_0.r15_2_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_2_ ),
    .Y(_02918_)
  );
  AOI22X1 _09553_ (
    .A( execution_unit_0.register_file_0.r6_2_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_2_ ),
    .Y(_02919_)
  );
  NAND2X1 _09554_ (
    .A(_02918_),
    .B(_02919_),
    .Y(_02920_)
  );
  AOI22X1 _09555_ (
    .A( execution_unit_0.register_file_0.r9_2_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_2_ ),
    .Y(_02921_)
  );
  AOI22X1 _09556_ (
    .A( execution_unit_0.alu_0.status_2_ ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_2_ ),
    .Y(_02922_)
  );
  NAND2X1 _09557_ (
    .A(_02921_),
    .B(_02922_),
    .Y(_02923_)
  );
  NOR2X1 _09558_ (
    .A(_02920_),
    .B(_02923_),
    .Y(_02924_)
  );
  NAND2X1 _09559_ (
    .A(_02917_),
    .B(_02924_),
    .Y( dbg_0.dbg_reg_din_2_ )
  );
  AOI22X1 _09560_ (
    .A( execution_unit_0.register_file_0.r1_3_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_3_ ),
    .Y(_02925_)
  );
  AOI22X1 _09561_ (
    .A( execution_unit_0.register_file_0.r5_3_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_3_ ),
    .Y(_02926_)
  );
  NAND2X1 _09562_ (
    .A(_02925_),
    .B(_02926_),
    .Y(_02927_)
  );
  AOI22X1 _09563_ (
    .A( execution_unit_0.register_file_0.r9_3_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_3_ ),
    .Y(_02928_)
  );
  AOI22X1 _09564_ (
    .A( execution_unit_0.gie ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.inst_dest_15_ ),
    .D( execution_unit_0.register_file_0.r15_3_ ),
    .Y(_02929_)
  );
  NAND2X1 _09565_ (
    .A(_02928_),
    .B(_02929_),
    .Y(_02930_)
  );
  NOR2X1 _09566_ (
    .A(_02927_),
    .B(_02930_),
    .Y(_02931_)
  );
  AOI22X1 _09567_ (
    .A( execution_unit_0.register_file_0.r7_3_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_6_ ),
    .D( execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02932_)
  );
  AOI22X1 _09568_ (
    .A( execution_unit_0.register_file_0.r12_3_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .C( dbg_0.UNUSED_pc_3_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02933_)
  );
  NAND2X1 _09569_ (
    .A(_02932_),
    .B(_02933_),
    .Y(_02934_)
  );
  AOI22X1 _09570_ (
    .A( execution_unit_0.register_file_0.r14_3_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_3_ ),
    .Y(_02935_)
  );
  AOI22X1 _09571_ (
    .A( execution_unit_0.register_file_0.r8_3_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_3_ ),
    .Y(_02936_)
  );
  NAND2X1 _09572_ (
    .A(_02935_),
    .B(_02936_),
    .Y(_02937_)
  );
  NOR2X1 _09573_ (
    .A(_02934_),
    .B(_02937_),
    .Y(_02938_)
  );
  NAND2X1 _09574_ (
    .A(_02931_),
    .B(_02938_),
    .Y( dbg_0.dbg_reg_din_3_ )
  );
  AOI22X1 _09575_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.register_file_0.r2_4_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_4_ ),
    .Y(_02939_)
  );
  AOI22X1 _09576_ (
    .A( execution_unit_0.register_file_0.r1_4_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02940_)
  );
  NAND2X1 _09577_ (
    .A(_02939_),
    .B(_02940_),
    .Y(_02941_)
  );
  AOI22X1 _09578_ (
    .A( execution_unit_0.register_file_0.r6_4_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02942_)
  );
  AOI22X1 _09579_ (
    .A( execution_unit_0.register_file_0.r14_4_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02943_)
  );
  NAND2X1 _09580_ (
    .A(_02942_),
    .B(_02943_),
    .Y(_02944_)
  );
  NOR2X1 _09581_ (
    .A(_02941_),
    .B(_02944_),
    .Y(_02945_)
  );
  AOI22X1 _09582_ (
    .A( execution_unit_0.register_file_0.r8_4_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_4_ ),
    .Y(_02946_)
  );
  AOI22X1 _09583_ (
    .A( execution_unit_0.register_file_0.r7_4_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_4_ ),
    .Y(_02947_)
  );
  NAND2X1 _09584_ (
    .A(_02946_),
    .B(_02947_),
    .Y(_02948_)
  );
  AOI22X1 _09585_ (
    .A( execution_unit_0.register_file_0.r15_4_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_4_ ),
    .Y(_02949_)
  );
  AOI22X1 _09586_ (
    .A( execution_unit_0.register_file_0.r9_4_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_4_ ),
    .Y(_02950_)
  );
  NAND2X1 _09587_ (
    .A(_02949_),
    .B(_02950_),
    .Y(_02951_)
  );
  NOR2X1 _09588_ (
    .A(_02948_),
    .B(_02951_),
    .Y(_02952_)
  );
  NAND2X1 _09589_ (
    .A(_02945_),
    .B(_02952_),
    .Y( dbg_0.dbg_reg_din_4_ )
  );
  AOI22X1 _09590_ (
    .A( execution_unit_0.register_file_0.r1_5_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_9_ ),
    .D( execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02953_)
  );
  AOI22X1 _09591_ (
    .A( clock_module_0.oscoff ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.inst_dest_7_ ),
    .D( execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02954_)
  );
  NAND2X1 _09592_ (
    .A(_02953_),
    .B(_02954_),
    .Y(_02955_)
  );
  AOI22X1 _09593_ (
    .A( execution_unit_0.register_file_0.r15_5_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_5_ ),
    .Y(_02956_)
  );
  AOI22X1 _09594_ (
    .A( execution_unit_0.register_file_0.r13_5_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_5_ ),
    .Y(_02957_)
  );
  NAND2X1 _09595_ (
    .A(_02956_),
    .B(_02957_),
    .Y(_02958_)
  );
  NOR2X1 _09596_ (
    .A(_02955_),
    .B(_02958_),
    .Y(_02959_)
  );
  AOI22X1 _09597_ (
    .A( execution_unit_0.register_file_0.r6_5_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_5_ ),
    .Y(_02960_)
  );
  AOI22X1 _09598_ (
    .A( execution_unit_0.register_file_0.r8_5_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_5_ ),
    .Y(_02961_)
  );
  NAND2X1 _09599_ (
    .A(_02960_),
    .B(_02961_),
    .Y(_02962_)
  );
  AOI22X1 _09600_ (
    .A( execution_unit_0.register_file_0.r5_5_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( dbg_0.UNUSED_pc_5_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02963_)
  );
  AOI22X1 _09601_ (
    .A( execution_unit_0.register_file_0.r4_5_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02964_)
  );
  NAND2X1 _09602_ (
    .A(_02963_),
    .B(_02964_),
    .Y(_02965_)
  );
  NOR2X1 _09603_ (
    .A(_02962_),
    .B(_02965_),
    .Y(_02966_)
  );
  NAND2X1 _09604_ (
    .A(_02959_),
    .B(_02966_),
    .Y( dbg_0.dbg_reg_din_5_ )
  );
  AOI22X1 _09605_ (
    .A( execution_unit_0.register_file_0.r7_6_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_6_ ),
    .Y(_02967_)
  );
  AOI22X1 _09606_ (
    .A( execution_unit_0.register_file_0.r15_6_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_6_ ),
    .Y(_02968_)
  );
  AND2X1 _09607_ (
    .A(_02967_),
    .B(_02968_),
    .Y(_02969_)
  );
  AOI22X1 _09608_ (
    .A( execution_unit_0.register_file_0.r8_6_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_6_ ),
    .Y(_02970_)
  );
  AOI22X1 _09609_ (
    .A( execution_unit_0.register_file_0.r1_6_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_6_ ),
    .Y(_02971_)
  );
  NAND3X1 _09610_ (
    .A(_02969_),
    .B(_02970_),
    .C(_02971_),
    .Y(_02972_)
  );
  AOI22X1 _09611_ (
    .A( execution_unit_0.register_file_0.r5_6_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_6_ ),
    .Y(_02973_)
  );
  INVX1 _09612_ (
    .A(_02973_),
    .Y(_02974_)
  );
  AOI21X1 _09613_ (
    .A( execution_unit_0.register_file_0.r11_6_ ),
    .B( execution_unit_0.inst_dest_11_ ),
    .C(_02974_),
    .Y(_02975_)
  );
  AOI22X1 _09614_ (
    .A( execution_unit_0.register_file_0.r6_6_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_6_ ),
    .Y(_02976_)
  );
  AOI22X1 _09615_ (
    .A( execution_unit_0.register_file_0.r9_6_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( dbg_0.UNUSED_pc_6_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02977_)
  );
  NAND3X1 _09616_ (
    .A(_02975_),
    .B(_02976_),
    .C(_02977_),
    .Y(_02978_)
  );
  OR2X1 _09617_ (
    .A(_02972_),
    .B(_02978_),
    .Y( dbg_0.dbg_reg_din_6_ )
  );
  AOI22X1 _09618_ (
    .A( execution_unit_0.register_file_0.r1_7_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_7_ ),
    .Y(_02979_)
  );
  AOI22X1 _09619_ (
    .A( execution_unit_0.register_file_0.r13_7_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_7_ ),
    .Y(_02980_)
  );
  NAND2X1 _09620_ (
    .A(_02979_),
    .B(_02980_),
    .Y(_02981_)
  );
  AOI22X1 _09621_ (
    .A( execution_unit_0.register_file_0.r9_7_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_7_ ),
    .Y(_02982_)
  );
  AOI22X1 _09622_ (
    .A( execution_unit_0.register_file_0.r15_7_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_7_ ),
    .Y(_02983_)
  );
  NAND2X1 _09623_ (
    .A(_02982_),
    .B(_02983_),
    .Y(_02984_)
  );
  NOR2X1 _09624_ (
    .A(_02981_),
    .B(_02984_),
    .Y(_02985_)
  );
  AOI22X1 _09625_ (
    .A( execution_unit_0.register_file_0.r7_7_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_6_ ),
    .D( execution_unit_0.register_file_0.r6_7_ ),
    .Y(_02986_)
  );
  AOI22X1 _09626_ (
    .A( execution_unit_0.register_file_0.r10_7_ ),
    .B( execution_unit_0.inst_dest_10_ ),
    .C( dbg_0.UNUSED_pc_7_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_02987_)
  );
  NAND2X1 _09627_ (
    .A(_02986_),
    .B(_02987_),
    .Y(_02988_)
  );
  AOI22X1 _09628_ (
    .A( clock_module_0.scg1 ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_7_ ),
    .Y(_02989_)
  );
  AOI22X1 _09629_ (
    .A( execution_unit_0.register_file_0.r8_7_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_7_ ),
    .Y(_02990_)
  );
  NAND2X1 _09630_ (
    .A(_02989_),
    .B(_02990_),
    .Y(_02991_)
  );
  NOR2X1 _09631_ (
    .A(_02988_),
    .B(_02991_),
    .Y(_02992_)
  );
  NAND2X1 _09632_ (
    .A(_02985_),
    .B(_02992_),
    .Y( dbg_0.dbg_reg_din_7_ )
  );
  AOI22X1 _09633_ (
    .A( execution_unit_0.register_file_0.r1_8_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_8_ ),
    .Y(_02993_)
  );
  AOI22X1 _09634_ (
    .A( execution_unit_0.register_file_0.r4_8_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_8_ ),
    .Y(_02994_)
  );
  NAND2X1 _09635_ (
    .A(_02993_),
    .B(_02994_),
    .Y(_02995_)
  );
  AOI22X1 _09636_ (
    .A( execution_unit_0.register_file_0.r8_8_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_8_ ),
    .Y(_02996_)
  );
  AOI22X1 _09637_ (
    .A( execution_unit_0.register_file_0.r15_8_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_8_ ),
    .Y(_02997_)
  );
  NAND2X1 _09638_ (
    .A(_02996_),
    .B(_02997_),
    .Y(_02998_)
  );
  NOR2X1 _09639_ (
    .A(_02995_),
    .B(_02998_),
    .Y(_02999_)
  );
  AOI22X1 _09640_ (
    .A( execution_unit_0.register_file_0.r7_8_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_6_ ),
    .D( execution_unit_0.register_file_0.r6_8_ ),
    .Y(_03000_)
  );
  AOI22X1 _09641_ (
    .A( execution_unit_0.register_file_0.r9_8_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_8_ ),
    .Y(_03001_)
  );
  NAND2X1 _09642_ (
    .A(_03000_),
    .B(_03001_),
    .Y(_03002_)
  );
  AOI22X1 _09643_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( dbg_0.UNUSED_pc_8_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03003_)
  );
  AOI22X1 _09644_ (
    .A( execution_unit_0.register_file_0.r13_8_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_8_ ),
    .Y(_03004_)
  );
  NAND2X1 _09645_ (
    .A(_03003_),
    .B(_03004_),
    .Y(_03005_)
  );
  NOR2X1 _09646_ (
    .A(_03002_),
    .B(_03005_),
    .Y(_03006_)
  );
  NAND2X1 _09647_ (
    .A(_02999_),
    .B(_03006_),
    .Y( dbg_0.dbg_reg_din_8_ )
  );
  NAND2X1 _09648_ (
    .A( execution_unit_0.register_file_0.r13_9_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_03007_)
  );
  NAND2X1 _09649_ (
    .A( execution_unit_0.register_file_0.r8_9_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .Y(_03008_)
  );
  AOI22X1 _09650_ (
    .A( execution_unit_0.register_file_0.r6_9_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( dbg_0.UNUSED_pc_9_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03009_)
  );
  AOI22X1 _09651_ (
    .A( execution_unit_0.register_file_0.r9_9_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_9_ ),
    .Y(_03010_)
  );
  AOI22X1 _09652_ (
    .A( execution_unit_0.register_file_0.r7_9_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_9_ ),
    .Y(_03011_)
  );
  AOI22X1 _09653_ (
    .A( execution_unit_0.register_file_0.r15_9_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_9_ ),
    .Y(_03012_)
  );
  AOI22X1 _09654_ (
    .A( execution_unit_0.register_file_0.r4_9_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_9_ ),
    .Y(_03013_)
  );
  NAND2X1 _09655_ (
    .A(_03012_),
    .B(_03013_),
    .Y(_03014_)
  );
  AOI21X1 _09656_ (
    .A( execution_unit_0.register_file_0.r11_9_ ),
    .B( execution_unit_0.inst_dest_11_ ),
    .C(_03014_),
    .Y(_03015_)
  );
  NAND3X1 _09657_ (
    .A(_03007_),
    .B(_03008_),
    .C(_03009_),
    .Y(_03016_)
  );
  AOI22X1 _09658_ (
    .A( execution_unit_0.register_file_0.r1_9_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_9_ ),
    .Y(_03017_)
  );
  NAND3X1 _09659_ (
    .A(_03010_),
    .B(_03011_),
    .C(_03017_),
    .Y(_03018_)
  );
  NOR2X1 _09660_ (
    .A(_03016_),
    .B(_03018_),
    .Y(_03019_)
  );
  NAND2X1 _09661_ (
    .A(_03015_),
    .B(_03019_),
    .Y( dbg_0.dbg_reg_din_9_ )
  );
  NAND2X1 _09662_ (
    .A( execution_unit_0.register_file_0.r3_10_ ),
    .B( execution_unit_0.inst_dest_3_ ),
    .Y(_03020_)
  );
  AOI22X1 _09663_ (
    .A( execution_unit_0.register_file_0.r1_10_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_10_ ),
    .Y(_03021_)
  );
  NAND2X1 _09664_ (
    .A(_03020_),
    .B(_03021_),
    .Y(_03022_)
  );
  AOI21X1 _09665_ (
    .A( execution_unit_0.register_file_0.r5_10_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C(_03022_),
    .Y(_03023_)
  );
  AOI22X1 _09666_ (
    .A( execution_unit_0.register_file_0.r8_10_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_10_ ),
    .Y(_03024_)
  );
  AOI22X1 _09667_ (
    .A( execution_unit_0.register_file_0.r6_10_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( dbg_0.UNUSED_pc_10_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03025_)
  );
  AND2X1 _09668_ (
    .A(_03024_),
    .B(_03025_),
    .Y(_03026_)
  );
  AOI22X1 _09669_ (
    .A( execution_unit_0.register_file_0.r7_10_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_15_ ),
    .D( execution_unit_0.register_file_0.r15_10_ ),
    .Y(_03027_)
  );
  AOI22X1 _09670_ (
    .A( execution_unit_0.register_file_0.r9_10_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_10_ ),
    .Y(_03028_)
  );
  AOI22X1 _09671_ (
    .A( execution_unit_0.register_file_0.r14_10_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_10_ ),
    .Y(_03029_)
  );
  NAND3X1 _09672_ (
    .A(_03027_),
    .B(_03028_),
    .C(_03029_),
    .Y(_03030_)
  );
  AOI21X1 _09673_ (
    .A( execution_unit_0.register_file_0.r10_10_ ),
    .B( execution_unit_0.inst_dest_10_ ),
    .C(_03030_),
    .Y(_03031_)
  );
  NAND3X1 _09674_ (
    .A(_03023_),
    .B(_03026_),
    .C(_03031_),
    .Y( dbg_0.dbg_reg_din_10_ )
  );
  NAND2X1 _09675_ (
    .A( execution_unit_0.register_file_0.r5_11_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .Y(_03032_)
  );
  NAND2X1 _09676_ (
    .A( execution_unit_0.register_file_0.r12_11_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_03033_)
  );
  AOI22X1 _09677_ (
    .A( execution_unit_0.register_file_0.r7_11_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_11_ ),
    .Y(_03034_)
  );
  AOI22X1 _09678_ (
    .A( execution_unit_0.register_file_0.r9_11_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( dbg_0.UNUSED_pc_11_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03035_)
  );
  NAND2X1 _09679_ (
    .A(_03033_),
    .B(_03035_),
    .Y(_03036_)
  );
  AOI21X1 _09680_ (
    .A( execution_unit_0.register_file_0.r1_11_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C(_03036_),
    .Y(_03037_)
  );
  AOI22X1 _09681_ (
    .A( execution_unit_0.register_file_0.r15_11_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_11_ ),
    .Y(_03038_)
  );
  AOI22X1 _09682_ (
    .A( execution_unit_0.register_file_0.r11_11_ ),
    .B( execution_unit_0.inst_dest_11_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_11_ ),
    .Y(_03039_)
  );
  NAND2X1 _09683_ (
    .A(_03038_),
    .B(_03039_),
    .Y(_03040_)
  );
  AOI21X1 _09684_ (
    .A( execution_unit_0.register_file_0.r13_11_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C(_03040_),
    .Y(_03041_)
  );
  AOI22X1 _09685_ (
    .A( execution_unit_0.register_file_0.r6_11_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_11_ ),
    .Y(_03042_)
  );
  NAND3X1 _09686_ (
    .A(_03032_),
    .B(_03034_),
    .C(_03042_),
    .Y(_03043_)
  );
  AOI21X1 _09687_ (
    .A( execution_unit_0.register_file_0.r8_11_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C(_03043_),
    .Y(_03044_)
  );
  NAND3X1 _09688_ (
    .A(_03037_),
    .B(_03041_),
    .C(_03044_),
    .Y( dbg_0.dbg_reg_din_11_ )
  );
  AOI22X1 _09689_ (
    .A( execution_unit_0.register_file_0.r12_12_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_12_ ),
    .Y(_03045_)
  );
  AOI22X1 _09690_ (
    .A( execution_unit_0.register_file_0.r8_12_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( dbg_0.UNUSED_pc_12_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03046_)
  );
  AND2X1 _09691_ (
    .A(_03045_),
    .B(_03046_),
    .Y(_03047_)
  );
  AOI22X1 _09692_ (
    .A( execution_unit_0.register_file_0.r7_12_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_12_ ),
    .Y(_03048_)
  );
  AOI22X1 _09693_ (
    .A( execution_unit_0.register_file_0.r9_12_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_12_ ),
    .Y(_03049_)
  );
  NAND3X1 _09694_ (
    .A(_03047_),
    .B(_03048_),
    .C(_03049_),
    .Y(_03050_)
  );
  AOI22X1 _09695_ (
    .A( execution_unit_0.register_file_0.r6_12_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_12_ ),
    .Y(_03051_)
  );
  INVX1 _09696_ (
    .A(_03051_),
    .Y(_03052_)
  );
  AOI21X1 _09697_ (
    .A( execution_unit_0.register_file_0.r14_12_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C(_03052_),
    .Y(_03053_)
  );
  AOI22X1 _09698_ (
    .A( execution_unit_0.register_file_0.r1_12_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_5_ ),
    .D( execution_unit_0.register_file_0.r5_12_ ),
    .Y(_03054_)
  );
  AOI22X1 _09699_ (
    .A( execution_unit_0.register_file_0.r15_12_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_12_ ),
    .Y(_03055_)
  );
  NAND3X1 _09700_ (
    .A(_03053_),
    .B(_03054_),
    .C(_03055_),
    .Y(_03056_)
  );
  OR2X1 _09701_ (
    .A(_03050_),
    .B(_03056_),
    .Y( dbg_0.dbg_reg_din_12_ )
  );
  AOI22X1 _09702_ (
    .A( execution_unit_0.register_file_0.r15_13_ ),
    .B( execution_unit_0.inst_dest_15_ ),
    .C( dbg_0.UNUSED_pc_13_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03057_)
  );
  AOI22X1 _09703_ (
    .A( execution_unit_0.register_file_0.r13_13_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_13_ ),
    .Y(_03058_)
  );
  AND2X1 _09704_ (
    .A(_03057_),
    .B(_03058_),
    .Y(_03059_)
  );
  AOI22X1 _09705_ (
    .A( execution_unit_0.register_file_0.r5_13_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( execution_unit_0.inst_dest_14_ ),
    .D( execution_unit_0.register_file_0.r14_13_ ),
    .Y(_03060_)
  );
  AOI22X1 _09706_ (
    .A( execution_unit_0.register_file_0.r8_13_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_7_ ),
    .D( execution_unit_0.register_file_0.r7_13_ ),
    .Y(_03061_)
  );
  NAND3X1 _09707_ (
    .A(_03059_),
    .B(_03060_),
    .C(_03061_),
    .Y(_03062_)
  );
  AOI22X1 _09708_ (
    .A( execution_unit_0.register_file_0.r1_13_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_13_ ),
    .Y(_03063_)
  );
  INVX1 _09709_ (
    .A(_03063_),
    .Y(_03064_)
  );
  AOI21X1 _09710_ (
    .A( execution_unit_0.register_file_0.r6_13_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C(_03064_),
    .Y(_03065_)
  );
  AOI22X1 _09711_ (
    .A( execution_unit_0.register_file_0.r4_13_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_13_ ),
    .Y(_03066_)
  );
  AOI22X1 _09712_ (
    .A( execution_unit_0.register_file_0.r9_13_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_13_ ),
    .Y(_03067_)
  );
  NAND3X1 _09713_ (
    .A(_03065_),
    .B(_03066_),
    .C(_03067_),
    .Y(_03068_)
  );
  OR2X1 _09714_ (
    .A(_03062_),
    .B(_03068_),
    .Y( dbg_0.dbg_reg_din_13_ )
  );
  AOI22X1 _09715_ (
    .A( execution_unit_0.register_file_0.r13_14_ ),
    .B( execution_unit_0.inst_dest_13_ ),
    .C( execution_unit_0.inst_dest_10_ ),
    .D( execution_unit_0.register_file_0.r10_14_ ),
    .Y(_03069_)
  );
  AOI22X1 _09716_ (
    .A( execution_unit_0.register_file_0.r4_14_ ),
    .B( execution_unit_0.inst_dest_4_ ),
    .C( dbg_0.UNUSED_pc_14_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03070_)
  );
  AND2X1 _09717_ (
    .A(_03069_),
    .B(_03070_),
    .Y(_03071_)
  );
  AOI22X1 _09718_ (
    .A( execution_unit_0.register_file_0.r9_14_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( execution_unit_0.inst_dest_15_ ),
    .D( execution_unit_0.register_file_0.r15_14_ ),
    .Y(_03072_)
  );
  AOI22X1 _09719_ (
    .A( execution_unit_0.register_file_0.r8_14_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_12_ ),
    .D( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_03073_)
  );
  NAND3X1 _09720_ (
    .A(_03071_),
    .B(_03072_),
    .C(_03073_),
    .Y(_03074_)
  );
  AOI22X1 _09721_ (
    .A( execution_unit_0.register_file_0.r14_14_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_14_ ),
    .Y(_03075_)
  );
  INVX1 _09722_ (
    .A(_03075_),
    .Y(_03076_)
  );
  AOI21X1 _09723_ (
    .A( execution_unit_0.register_file_0.r7_14_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C(_03076_),
    .Y(_03077_)
  );
  AOI22X1 _09724_ (
    .A( execution_unit_0.register_file_0.r1_14_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .C( execution_unit_0.inst_dest_6_ ),
    .D( execution_unit_0.register_file_0.r6_14_ ),
    .Y(_03078_)
  );
  AOI22X1 _09725_ (
    .A( execution_unit_0.register_file_0.r5_14_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_14_ ),
    .Y(_03079_)
  );
  NAND3X1 _09726_ (
    .A(_03077_),
    .B(_03078_),
    .C(_03079_),
    .Y(_03080_)
  );
  OR2X1 _09727_ (
    .A(_03074_),
    .B(_03080_),
    .Y( dbg_0.dbg_reg_din_14_ )
  );
  NAND2X1 _09728_ (
    .A( execution_unit_0.register_file_0.r1_15_ ),
    .B( execution_unit_0.inst_dest_1_ ),
    .Y(_03081_)
  );
  NAND2X1 _09729_ (
    .A( execution_unit_0.register_file_0.r12_15_ ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_03082_)
  );
  AOI22X1 _09730_ (
    .A( execution_unit_0.register_file_0.r9_15_ ),
    .B( execution_unit_0.inst_dest_9_ ),
    .C( dbg_0.UNUSED_pc_15_ ),
    .D( execution_unit_0.inst_dest_0_ ),
    .Y(_03083_)
  );
  NAND2X1 _09731_ (
    .A(_03082_),
    .B(_03083_),
    .Y(_03084_)
  );
  AOI22X1 _09732_ (
    .A( execution_unit_0.register_file_0.r10_15_ ),
    .B( execution_unit_0.inst_dest_10_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_15_ ),
    .Y(_03085_)
  );
  AOI22X1 _09733_ (
    .A( execution_unit_0.register_file_0.r5_15_ ),
    .B( execution_unit_0.inst_dest_5_ ),
    .C( execution_unit_0.inst_dest_4_ ),
    .D( execution_unit_0.register_file_0.r4_15_ ),
    .Y(_03086_)
  );
  NAND3X1 _09734_ (
    .A(_03081_),
    .B(_03085_),
    .C(_03086_),
    .Y(_03087_)
  );
  NOR2X1 _09735_ (
    .A(_03084_),
    .B(_03087_),
    .Y(_03088_)
  );
  AOI22X1 _09736_ (
    .A( execution_unit_0.register_file_0.r7_15_ ),
    .B( execution_unit_0.inst_dest_7_ ),
    .C( execution_unit_0.inst_dest_11_ ),
    .D( execution_unit_0.register_file_0.r11_15_ ),
    .Y(_03089_)
  );
  AOI22X1 _09737_ (
    .A( execution_unit_0.register_file_0.r8_15_ ),
    .B( execution_unit_0.inst_dest_8_ ),
    .C( execution_unit_0.inst_dest_13_ ),
    .D( execution_unit_0.register_file_0.r13_15_ ),
    .Y(_03090_)
  );
  AOI22X1 _09738_ (
    .A( execution_unit_0.register_file_0.r6_15_ ),
    .B( execution_unit_0.inst_dest_6_ ),
    .C( execution_unit_0.inst_dest_15_ ),
    .D( execution_unit_0.register_file_0.r15_15_ ),
    .Y(_03091_)
  );
  NAND3X1 _09739_ (
    .A(_03089_),
    .B(_03090_),
    .C(_03091_),
    .Y(_03092_)
  );
  AOI21X1 _09740_ (
    .A( execution_unit_0.register_file_0.r14_15_ ),
    .B( execution_unit_0.inst_dest_14_ ),
    .C(_03092_),
    .Y(_03093_)
  );
  NAND2X1 _09741_ (
    .A(_03088_),
    .B(_03093_),
    .Y( dbg_0.dbg_reg_din_15_ )
  );
  INVX1 _09742_ (
    .A(_06327_),
    .Y(_01902_)
  );
  INVX1 _09743_ (
    .A(_06327_),
    .Y(_01903_)
  );
  INVX1 _09744_ (
    .A(_06327_),
    .Y(_01904_)
  );
  INVX1 _09745_ (
    .A(_06327_),
    .Y(_01905_)
  );
  INVX1 _09746_ (
    .A(_06327_),
    .Y(_01906_)
  );
  INVX1 _09747_ (
    .A(_06327_),
    .Y(_01907_)
  );
  INVX1 _09748_ (
    .A(_06327_),
    .Y(_01908_)
  );
  INVX1 _09749_ (
    .A(_06327_),
    .Y(_01909_)
  );
  INVX1 _09750_ (
    .A(_06327_),
    .Y(_01910_)
  );
  INVX1 _09751_ (
    .A(_06327_),
    .Y(_01911_)
  );
  INVX1 _09752_ (
    .A(_06327_),
    .Y(_01912_)
  );
  INVX1 _09753_ (
    .A(_06327_),
    .Y(_01913_)
  );
  INVX1 _09754_ (
    .A(_06327_),
    .Y(_01914_)
  );
  INVX1 _09755_ (
    .A(_06327_),
    .Y(_01915_)
  );
  INVX1 _09756_ (
    .A(_06327_),
    .Y(_01916_)
  );
  INVX1 _09757_ (
    .A(_06327_),
    .Y(_01917_)
  );
  INVX1 _09758_ (
    .A(_06327_),
    .Y(_01918_)
  );
  INVX1 _09759_ (
    .A(_06327_),
    .Y(_01919_)
  );
  INVX1 _09760_ (
    .A(_06327_),
    .Y(_01920_)
  );
  INVX1 _09761_ (
    .A(_06327_),
    .Y(_01921_)
  );
  INVX1 _09762_ (
    .A(_06327_),
    .Y(_01922_)
  );
  INVX1 _09763_ (
    .A(_06327_),
    .Y(_01923_)
  );
  INVX1 _09764_ (
    .A(_06327_),
    .Y(_01924_)
  );
  INVX1 _09765_ (
    .A(_06327_),
    .Y(_01925_)
  );
  INVX1 _09766_ (
    .A(_06327_),
    .Y(_01926_)
  );
  INVX1 _09767_ (
    .A(_06327_),
    .Y(_01927_)
  );
  INVX1 _09768_ (
    .A(_06327_),
    .Y(_01928_)
  );
  INVX1 _09769_ (
    .A(_06327_),
    .Y(_01929_)
  );
  INVX1 _09770_ (
    .A(_06327_),
    .Y(_01930_)
  );
  INVX1 _09771_ (
    .A(_06327_),
    .Y(_01931_)
  );
  INVX1 _09772_ (
    .A(_06327_),
    .Y(_01932_)
  );
  INVX1 _09773_ (
    .A(_06327_),
    .Y(_01933_)
  );
  INVX1 _09774_ (
    .A(_06327_),
    .Y(_01934_)
  );
  INVX1 _09775_ (
    .A(_06327_),
    .Y(_01935_)
  );
  INVX1 _09776_ (
    .A(_06327_),
    .Y(_01936_)
  );
  INVX1 _09777_ (
    .A(_06327_),
    .Y(_01937_)
  );
  INVX1 _09778_ (
    .A(_06327_),
    .Y(_01938_)
  );
  INVX1 _09779_ (
    .A(_06327_),
    .Y(_01939_)
  );
  INVX1 _09780_ (
    .A(_06327_),
    .Y(_01940_)
  );
  INVX1 _09781_ (
    .A(_06327_),
    .Y(_01941_)
  );
  INVX1 _09782_ (
    .A(_06327_),
    .Y(_01942_)
  );
  INVX1 _09783_ (
    .A(_06327_),
    .Y(_01943_)
  );
  INVX1 _09784_ (
    .A(_06327_),
    .Y(_01944_)
  );
  INVX1 _09785_ (
    .A(_06327_),
    .Y(_01945_)
  );
  INVX1 _09786_ (
    .A(_06327_),
    .Y(_01946_)
  );
  INVX1 _09787_ (
    .A(_06327_),
    .Y(_01947_)
  );
  INVX1 _09788_ (
    .A(_06327_),
    .Y(_01948_)
  );
  INVX1 _09789_ (
    .A(_06327_),
    .Y(_01949_)
  );
  INVX1 _09790_ (
    .A(_06327_),
    .Y(_01950_)
  );
  INVX1 _09791_ (
    .A(_06327_),
    .Y(_01951_)
  );
  INVX1 _09792_ (
    .A(_06327_),
    .Y(_01952_)
  );
  INVX1 _09793_ (
    .A(_06327_),
    .Y(_01953_)
  );
  INVX1 _09794_ (
    .A(_06327_),
    .Y(_01954_)
  );
  INVX1 _09795_ (
    .A(_06327_),
    .Y(_01955_)
  );
  INVX1 _09796_ (
    .A(_06327_),
    .Y(_01956_)
  );
  INVX1 _09797_ (
    .A(_06327_),
    .Y(_01957_)
  );
  INVX1 _09798_ (
    .A(_06327_),
    .Y(_01958_)
  );
  INVX1 _09799_ (
    .A(_06327_),
    .Y(_01959_)
  );
  INVX1 _09800_ (
    .A(_06327_),
    .Y(_01960_)
  );
  INVX1 _09801_ (
    .A(_06327_),
    .Y(_01961_)
  );
  INVX1 _09802_ (
    .A(_06327_),
    .Y(_01962_)
  );
  INVX1 _09803_ (
    .A(_06327_),
    .Y(_01963_)
  );
  INVX1 _09804_ (
    .A(_06327_),
    .Y(_01964_)
  );
  INVX1 _09805_ (
    .A(_06327_),
    .Y(_01965_)
  );
  INVX1 _09806_ (
    .A(_06327_),
    .Y(_01966_)
  );
  INVX1 _09807_ (
    .A(_06327_),
    .Y(_01967_)
  );
  INVX1 _09808_ (
    .A(_06327_),
    .Y(_01968_)
  );
  INVX1 _09809_ (
    .A(_06327_),
    .Y(_01969_)
  );
  INVX1 _09810_ (
    .A(_06327_),
    .Y(_01970_)
  );
  INVX1 _09811_ (
    .A(_06327_),
    .Y(_01971_)
  );
  INVX1 _09812_ (
    .A(_06327_),
    .Y(_01972_)
  );
  INVX1 _09813_ (
    .A(_06327_),
    .Y(_01973_)
  );
  INVX1 _09814_ (
    .A(_06327_),
    .Y(_01974_)
  );
  INVX1 _09815_ (
    .A(_06327_),
    .Y(_01975_)
  );
  INVX1 _09816_ (
    .A(_06327_),
    .Y(_01976_)
  );
  INVX1 _09817_ (
    .A(_06327_),
    .Y(_01977_)
  );
  INVX1 _09818_ (
    .A(_06327_),
    .Y(_01978_)
  );
  INVX1 _09819_ (
    .A(_06327_),
    .Y(_01979_)
  );
  INVX1 _09820_ (
    .A(_06327_),
    .Y(_01980_)
  );
  INVX1 _09821_ (
    .A(_06327_),
    .Y(_01981_)
  );
  INVX1 _09822_ (
    .A(_06327_),
    .Y(_01982_)
  );
  INVX1 _09823_ (
    .A(_06327_),
    .Y(_01983_)
  );
  INVX1 _09824_ (
    .A(_06327_),
    .Y(_01984_)
  );
  INVX1 _09825_ (
    .A(_06327_),
    .Y(_01985_)
  );
  INVX1 _09826_ (
    .A(_06327_),
    .Y(_01986_)
  );
  INVX1 _09827_ (
    .A(_06327_),
    .Y(_01987_)
  );
  INVX1 _09828_ (
    .A(_06327_),
    .Y(_01988_)
  );
  INVX1 _09829_ (
    .A(_06327_),
    .Y(_01989_)
  );
  INVX1 _09830_ (
    .A(_06327_),
    .Y(_01990_)
  );
  INVX1 _09831_ (
    .A(_06327_),
    .Y(_01991_)
  );
  INVX1 _09832_ (
    .A(_06327_),
    .Y(_01992_)
  );
  INVX1 _09833_ (
    .A(_06327_),
    .Y(_01993_)
  );
  INVX1 _09834_ (
    .A(_06327_),
    .Y(_01994_)
  );
  INVX1 _09835_ (
    .A(_06327_),
    .Y(_01995_)
  );
  INVX1 _09836_ (
    .A(_06327_),
    .Y(_01996_)
  );
  INVX1 _09837_ (
    .A(_06327_),
    .Y(_01997_)
  );
  INVX1 _09838_ (
    .A(_06327_),
    .Y(_01998_)
  );
  INVX1 _09839_ (
    .A(_06327_),
    .Y(_01999_)
  );
  INVX1 _09840_ (
    .A(_06327_),
    .Y(_02000_)
  );
  INVX1 _09841_ (
    .A(_06327_),
    .Y(_02001_)
  );
  INVX1 _09842_ (
    .A(_06327_),
    .Y(_02002_)
  );
  INVX1 _09843_ (
    .A(_06327_),
    .Y(_02003_)
  );
  INVX1 _09844_ (
    .A(_06327_),
    .Y(_02004_)
  );
  INVX1 _09845_ (
    .A(_06327_),
    .Y(_02005_)
  );
  INVX1 _09846_ (
    .A(_06327_),
    .Y(_02006_)
  );
  INVX1 _09847_ (
    .A(_06327_),
    .Y(_02007_)
  );
  INVX1 _09848_ (
    .A(_06327_),
    .Y(_02008_)
  );
  INVX1 _09849_ (
    .A(_06327_),
    .Y(_02009_)
  );
  INVX1 _09850_ (
    .A(_06327_),
    .Y(_02010_)
  );
  INVX1 _09851_ (
    .A(_06327_),
    .Y(_02011_)
  );
  INVX1 _09852_ (
    .A(_06327_),
    .Y(_02012_)
  );
  INVX1 _09853_ (
    .A(_06327_),
    .Y(_02013_)
  );
  INVX1 _09854_ (
    .A(_06327_),
    .Y(_02014_)
  );
  INVX1 _09855_ (
    .A(_06327_),
    .Y(_02015_)
  );
  INVX1 _09856_ (
    .A(_06327_),
    .Y(_02016_)
  );
  INVX1 _09857_ (
    .A(_06327_),
    .Y(_02017_)
  );
  INVX1 _09858_ (
    .A(_06327_),
    .Y(_02018_)
  );
  INVX1 _09859_ (
    .A(_06327_),
    .Y(_02019_)
  );
  INVX1 _09860_ (
    .A(_06327_),
    .Y(_02020_)
  );
  INVX1 _09861_ (
    .A(_06327_),
    .Y(_02021_)
  );
  INVX1 _09862_ (
    .A(_06327_),
    .Y(_02022_)
  );
  INVX1 _09863_ (
    .A(_06327_),
    .Y(_02023_)
  );
  INVX1 _09864_ (
    .A(_06327_),
    .Y(_02024_)
  );
  INVX1 _09865_ (
    .A(_06327_),
    .Y(_02025_)
  );
  INVX1 _09866_ (
    .A(_06327_),
    .Y(_02026_)
  );
  INVX1 _09867_ (
    .A(_06327_),
    .Y(_02027_)
  );
  INVX1 _09868_ (
    .A(_06327_),
    .Y(_02028_)
  );
  INVX1 _09869_ (
    .A(_06327_),
    .Y(_02029_)
  );
  INVX1 _09870_ (
    .A(_06327_),
    .Y(_02030_)
  );
  INVX1 _09871_ (
    .A(_06327_),
    .Y(_02031_)
  );
  INVX1 _09872_ (
    .A(_06327_),
    .Y(_02032_)
  );
  INVX1 _09873_ (
    .A(_06327_),
    .Y(_02033_)
  );
  INVX1 _09874_ (
    .A(_06327_),
    .Y(_02034_)
  );
  INVX1 _09875_ (
    .A(_06327_),
    .Y(_02035_)
  );
  INVX1 _09876_ (
    .A(_06327_),
    .Y(_02036_)
  );
  INVX1 _09877_ (
    .A(_06327_),
    .Y(_02037_)
  );
  INVX1 _09878_ (
    .A(_06327_),
    .Y(_02038_)
  );
  INVX1 _09879_ (
    .A(_06327_),
    .Y(_02039_)
  );
  INVX1 _09880_ (
    .A(_06327_),
    .Y(_02040_)
  );
  INVX1 _09881_ (
    .A(_06327_),
    .Y(_02041_)
  );
  INVX1 _09882_ (
    .A(_06327_),
    .Y(_02042_)
  );
  INVX1 _09883_ (
    .A(_06327_),
    .Y(_02043_)
  );
  INVX1 _09884_ (
    .A(_06327_),
    .Y(_02044_)
  );
  INVX1 _09885_ (
    .A(_06327_),
    .Y(_02045_)
  );
  INVX1 _09886_ (
    .A(_06327_),
    .Y(_02046_)
  );
  INVX1 _09887_ (
    .A(_06327_),
    .Y(_02047_)
  );
  INVX1 _09888_ (
    .A(_06327_),
    .Y(_02048_)
  );
  INVX1 _09889_ (
    .A(_06327_),
    .Y(_02049_)
  );
  INVX1 _09890_ (
    .A(_06327_),
    .Y(_02050_)
  );
  INVX1 _09891_ (
    .A(_06327_),
    .Y(_02051_)
  );
  INVX1 _09892_ (
    .A(_06327_),
    .Y(_02052_)
  );
  INVX1 _09893_ (
    .A(_06327_),
    .Y(_02053_)
  );
  INVX1 _09894_ (
    .A(_06327_),
    .Y(_02054_)
  );
  INVX1 _09895_ (
    .A(_06327_),
    .Y(_02055_)
  );
  INVX1 _09896_ (
    .A(_06327_),
    .Y(_02056_)
  );
  INVX1 _09897_ (
    .A(_06327_),
    .Y(_02057_)
  );
  INVX1 _09898_ (
    .A(_06327_),
    .Y(_02058_)
  );
  INVX1 _09899_ (
    .A(_06327_),
    .Y(_02059_)
  );
  INVX1 _09900_ (
    .A(_06327_),
    .Y(_02060_)
  );
  INVX1 _09901_ (
    .A(_06327_),
    .Y(_02061_)
  );
  INVX1 _09902_ (
    .A(_06327_),
    .Y(_02062_)
  );
  INVX1 _09903_ (
    .A(_06327_),
    .Y(_02063_)
  );
  INVX1 _09904_ (
    .A(_06327_),
    .Y(_02064_)
  );
  INVX1 _09905_ (
    .A(_06327_),
    .Y(_02065_)
  );
  INVX1 _09906_ (
    .A(_06327_),
    .Y(_02066_)
  );
  INVX1 _09907_ (
    .A(_06327_),
    .Y(_02067_)
  );
  INVX1 _09908_ (
    .A(_06327_),
    .Y(_02068_)
  );
  INVX1 _09909_ (
    .A(_06327_),
    .Y(_02069_)
  );
  INVX1 _09910_ (
    .A(_06327_),
    .Y(_02070_)
  );
  INVX1 _09911_ (
    .A(_06327_),
    .Y(_02071_)
  );
  INVX1 _09912_ (
    .A(_06327_),
    .Y(_02072_)
  );
  INVX1 _09913_ (
    .A(_06327_),
    .Y(_02073_)
  );
  INVX1 _09914_ (
    .A(_06327_),
    .Y(_02074_)
  );
  INVX1 _09915_ (
    .A(_06327_),
    .Y(_02075_)
  );
  INVX1 _09916_ (
    .A(_06327_),
    .Y(_02076_)
  );
  INVX1 _09917_ (
    .A(_06327_),
    .Y(_02077_)
  );
  INVX1 _09918_ (
    .A(_06327_),
    .Y(_02078_)
  );
  INVX1 _09919_ (
    .A(_06327_),
    .Y(_02079_)
  );
  INVX1 _09920_ (
    .A(_06327_),
    .Y(_02080_)
  );
  INVX1 _09921_ (
    .A(_06327_),
    .Y(_02081_)
  );
  INVX1 _09922_ (
    .A(_06327_),
    .Y(_02082_)
  );
  INVX1 _09923_ (
    .A(_06327_),
    .Y(_02083_)
  );
  INVX1 _09924_ (
    .A(_06327_),
    .Y(_02084_)
  );
  INVX1 _09925_ (
    .A(_06327_),
    .Y(_02085_)
  );
  INVX1 _09926_ (
    .A(_06327_),
    .Y(_02086_)
  );
  INVX1 _09927_ (
    .A(_06327_),
    .Y(_02087_)
  );
  INVX1 _09928_ (
    .A(_06327_),
    .Y(_02088_)
  );
  INVX1 _09929_ (
    .A(_06327_),
    .Y(_02089_)
  );
  INVX1 _09930_ (
    .A(_06327_),
    .Y(_02090_)
  );
  INVX1 _09931_ (
    .A(_06327_),
    .Y(_02091_)
  );
  INVX1 _09932_ (
    .A(_06327_),
    .Y(_02092_)
  );
  INVX1 _09933_ (
    .A(_06327_),
    .Y(_02093_)
  );
  INVX1 _09934_ (
    .A(_06327_),
    .Y(_02094_)
  );
  INVX1 _09935_ (
    .A(_06327_),
    .Y(_02095_)
  );
  INVX1 _09936_ (
    .A(_06327_),
    .Y(_02096_)
  );
  INVX1 _09937_ (
    .A(_06327_),
    .Y(_02097_)
  );
  INVX1 _09938_ (
    .A(_06327_),
    .Y(_02098_)
  );
  INVX1 _09939_ (
    .A(_06327_),
    .Y(_02099_)
  );
  INVX1 _09940_ (
    .A(_06327_),
    .Y(_02100_)
  );
  INVX1 _09941_ (
    .A(_06327_),
    .Y(_02101_)
  );
  INVX1 _09942_ (
    .A(_06327_),
    .Y(_02102_)
  );
  INVX1 _09943_ (
    .A(_06327_),
    .Y(_02103_)
  );
  INVX1 _09944_ (
    .A(_06327_),
    .Y(_02104_)
  );
  INVX1 _09945_ (
    .A(_06327_),
    .Y(_02105_)
  );
  INVX1 _09946_ (
    .A(_06327_),
    .Y(_02106_)
  );
  INVX1 _09947_ (
    .A(_06327_),
    .Y(_02107_)
  );
  INVX1 _09948_ (
    .A(_06327_),
    .Y(_02108_)
  );
  INVX1 _09949_ (
    .A(_06327_),
    .Y(_02109_)
  );
  INVX1 _09950_ (
    .A(_06327_),
    .Y(_02110_)
  );
  INVX1 _09951_ (
    .A(_06327_),
    .Y(_02111_)
  );
  INVX1 _09952_ (
    .A(_06327_),
    .Y(_02112_)
  );
  INVX1 _09953_ (
    .A(_06327_),
    .Y(_02113_)
  );
  INVX1 _09954_ (
    .A(_06327_),
    .Y(_02114_)
  );
  INVX1 _09955_ (
    .A(_06327_),
    .Y(_02115_)
  );
  INVX1 _09956_ (
    .A(_06327_),
    .Y(_02116_)
  );
  INVX1 _09957_ (
    .A(_06327_),
    .Y(_02117_)
  );
  INVX1 _09958_ (
    .A(_06327_),
    .Y(_02118_)
  );
  INVX1 _09959_ (
    .A(_06327_),
    .Y(_02119_)
  );
  INVX1 _09960_ (
    .A(_06327_),
    .Y(_02120_)
  );
  INVX1 _09961_ (
    .A(_06327_),
    .Y(_02121_)
  );
  INVX1 _09962_ (
    .A(_06327_),
    .Y(_02122_)
  );
  INVX1 _09963_ (
    .A(_06327_),
    .Y(_02123_)
  );
  INVX1 _09964_ (
    .A(_06327_),
    .Y(_02124_)
  );
  INVX1 _09965_ (
    .A(_06327_),
    .Y(_02125_)
  );
  INVX1 _09966_ (
    .A(_06327_),
    .Y(_02126_)
  );
  INVX1 _09967_ (
    .A(_06327_),
    .Y(_02127_)
  );
  INVX1 _09968_ (
    .A(_06327_),
    .Y(_02128_)
  );
  INVX1 _09969_ (
    .A(_06327_),
    .Y(_02129_)
  );
  INVX1 _09970_ (
    .A(_06327_),
    .Y(_02130_)
  );
  INVX1 _09971_ (
    .A(_06327_),
    .Y(_02131_)
  );
  DFFSR _09972_ (
    .CLK(dco_clk),
    .D(_02132_),
    .Q( execution_unit_0.alu_0.status_1_ ),
    .R(_01901_),
    .S(1'h1)
  );
  DFFSR _09973_ (
    .CLK(dco_clk),
    .D(_02133_),
    .Q( execution_unit_0.alu_0.status_2_ ),
    .R(_01902_),
    .S(1'h1)
  );
  DFFSR _09974_ (
    .CLK(dco_clk),
    .D(_02134_),
    .Q( execution_unit_0.gie ),
    .R(_01903_),
    .S(1'h1)
  );
  DFFSR _09975_ (
    .CLK(dco_clk),
    .D(_02135_),
    .Q( clock_module_0.oscoff ),
    .R(_01904_),
    .S(1'h1)
  );
  DFFSR _09976_ (
    .CLK(dco_clk),
    .D(_02136_),
    .Q( clock_module_0.scg1 ),
    .R(_01905_),
    .S(1'h1)
  );
  DFFSR _09977_ (
    .CLK(dco_clk),
    .D(_02137_),
    .Q( execution_unit_0.alu_0.status_3_ ),
    .R(_01906_),
    .S(1'h1)
  );
  DFFSR _09978_ (
    .CLK(dco_clk),
    .D(_02138_),
    .Q( execution_unit_0.register_file_0.r15_0_ ),
    .R(_01907_),
    .S(1'h1)
  );
  DFFSR _09979_ (
    .CLK(dco_clk),
    .D(_02139_),
    .Q( execution_unit_0.register_file_0.r15_1_ ),
    .R(_01908_),
    .S(1'h1)
  );
  DFFSR _09980_ (
    .CLK(dco_clk),
    .D(_02140_),
    .Q( execution_unit_0.register_file_0.r15_2_ ),
    .R(_01909_),
    .S(1'h1)
  );
  DFFSR _09981_ (
    .CLK(dco_clk),
    .D(_02141_),
    .Q( execution_unit_0.register_file_0.r15_3_ ),
    .R(_01910_),
    .S(1'h1)
  );
  DFFSR _09982_ (
    .CLK(dco_clk),
    .D(_02142_),
    .Q( execution_unit_0.register_file_0.r15_4_ ),
    .R(_01911_),
    .S(1'h1)
  );
  DFFSR _09983_ (
    .CLK(dco_clk),
    .D(_02143_),
    .Q( execution_unit_0.register_file_0.r15_5_ ),
    .R(_01912_),
    .S(1'h1)
  );
  DFFSR _09984_ (
    .CLK(dco_clk),
    .D(_02144_),
    .Q( execution_unit_0.register_file_0.r15_6_ ),
    .R(_01913_),
    .S(1'h1)
  );
  DFFSR _09985_ (
    .CLK(dco_clk),
    .D(_02145_),
    .Q( execution_unit_0.register_file_0.r15_7_ ),
    .R(_01914_),
    .S(1'h1)
  );
  DFFSR _09986_ (
    .CLK(dco_clk),
    .D(_02146_),
    .Q( execution_unit_0.register_file_0.r15_8_ ),
    .R(_01915_),
    .S(1'h1)
  );
  DFFSR _09987_ (
    .CLK(dco_clk),
    .D(_02147_),
    .Q( execution_unit_0.register_file_0.r15_9_ ),
    .R(_01916_),
    .S(1'h1)
  );
  DFFSR _09988_ (
    .CLK(dco_clk),
    .D(_02148_),
    .Q( execution_unit_0.register_file_0.r15_10_ ),
    .R(_01917_),
    .S(1'h1)
  );
  DFFSR _09989_ (
    .CLK(dco_clk),
    .D(_02149_),
    .Q( execution_unit_0.register_file_0.r15_11_ ),
    .R(_01918_),
    .S(1'h1)
  );
  DFFSR _09990_ (
    .CLK(dco_clk),
    .D(_02150_),
    .Q( execution_unit_0.register_file_0.r15_12_ ),
    .R(_01919_),
    .S(1'h1)
  );
  DFFSR _09991_ (
    .CLK(dco_clk),
    .D(_02151_),
    .Q( execution_unit_0.register_file_0.r15_13_ ),
    .R(_01920_),
    .S(1'h1)
  );
  DFFSR _09992_ (
    .CLK(dco_clk),
    .D(_02152_),
    .Q( execution_unit_0.register_file_0.r15_14_ ),
    .R(_01921_),
    .S(1'h1)
  );
  DFFSR _09993_ (
    .CLK(dco_clk),
    .D(_02153_),
    .Q( execution_unit_0.register_file_0.r15_15_ ),
    .R(_01922_),
    .S(1'h1)
  );
  DFFSR _09994_ (
    .CLK(dco_clk),
    .D(_02154_),
    .Q( execution_unit_0.register_file_0.r14_0_ ),
    .R(_01923_),
    .S(1'h1)
  );
  DFFSR _09995_ (
    .CLK(dco_clk),
    .D(_02155_),
    .Q( execution_unit_0.register_file_0.r14_1_ ),
    .R(_01924_),
    .S(1'h1)
  );
  DFFSR _09996_ (
    .CLK(dco_clk),
    .D(_02156_),
    .Q( execution_unit_0.register_file_0.r14_2_ ),
    .R(_01925_),
    .S(1'h1)
  );
  DFFSR _09997_ (
    .CLK(dco_clk),
    .D(_02157_),
    .Q( execution_unit_0.register_file_0.r14_3_ ),
    .R(_01926_),
    .S(1'h1)
  );
  DFFSR _09998_ (
    .CLK(dco_clk),
    .D(_02158_),
    .Q( execution_unit_0.register_file_0.r14_4_ ),
    .R(_01927_),
    .S(1'h1)
  );
  DFFSR _09999_ (
    .CLK(dco_clk),
    .D(_02159_),
    .Q( execution_unit_0.register_file_0.r14_5_ ),
    .R(_01928_),
    .S(1'h1)
  );
  DFFSR _10000_ (
    .CLK(dco_clk),
    .D(_02160_),
    .Q( execution_unit_0.register_file_0.r14_6_ ),
    .R(_01929_),
    .S(1'h1)
  );
  DFFSR _10001_ (
    .CLK(dco_clk),
    .D(_02161_),
    .Q( execution_unit_0.register_file_0.r14_7_ ),
    .R(_01930_),
    .S(1'h1)
  );
  DFFSR _10002_ (
    .CLK(dco_clk),
    .D(_02162_),
    .Q( execution_unit_0.register_file_0.r14_8_ ),
    .R(_01931_),
    .S(1'h1)
  );
  DFFSR _10003_ (
    .CLK(dco_clk),
    .D(_02163_),
    .Q( execution_unit_0.register_file_0.r14_9_ ),
    .R(_01932_),
    .S(1'h1)
  );
  DFFSR _10004_ (
    .CLK(dco_clk),
    .D(_02164_),
    .Q( execution_unit_0.register_file_0.r14_10_ ),
    .R(_01933_),
    .S(1'h1)
  );
  DFFSR _10005_ (
    .CLK(dco_clk),
    .D(_02165_),
    .Q( execution_unit_0.register_file_0.r14_11_ ),
    .R(_01934_),
    .S(1'h1)
  );
  DFFSR _10006_ (
    .CLK(dco_clk),
    .D(_02166_),
    .Q( execution_unit_0.register_file_0.r14_12_ ),
    .R(_01935_),
    .S(1'h1)
  );
  DFFSR _10007_ (
    .CLK(dco_clk),
    .D(_02167_),
    .Q( execution_unit_0.register_file_0.r14_13_ ),
    .R(_01936_),
    .S(1'h1)
  );
  DFFSR _10008_ (
    .CLK(dco_clk),
    .D(_02168_),
    .Q( execution_unit_0.register_file_0.r14_14_ ),
    .R(_01937_),
    .S(1'h1)
  );
  DFFSR _10009_ (
    .CLK(dco_clk),
    .D(_02169_),
    .Q( execution_unit_0.register_file_0.r14_15_ ),
    .R(_01938_),
    .S(1'h1)
  );
  DFFSR _10010_ (
    .CLK(dco_clk),
    .D(_02170_),
    .Q( execution_unit_0.register_file_0.r13_0_ ),
    .R(_01939_),
    .S(1'h1)
  );
  DFFSR _10011_ (
    .CLK(dco_clk),
    .D(_02171_),
    .Q( execution_unit_0.register_file_0.r13_1_ ),
    .R(_01940_),
    .S(1'h1)
  );
  DFFSR _10012_ (
    .CLK(dco_clk),
    .D(_02172_),
    .Q( execution_unit_0.register_file_0.r13_2_ ),
    .R(_01941_),
    .S(1'h1)
  );
  DFFSR _10013_ (
    .CLK(dco_clk),
    .D(_02173_),
    .Q( execution_unit_0.register_file_0.r13_3_ ),
    .R(_01942_),
    .S(1'h1)
  );
  DFFSR _10014_ (
    .CLK(dco_clk),
    .D(_02174_),
    .Q( execution_unit_0.register_file_0.r13_4_ ),
    .R(_01943_),
    .S(1'h1)
  );
  DFFSR _10015_ (
    .CLK(dco_clk),
    .D(_02175_),
    .Q( execution_unit_0.register_file_0.r13_5_ ),
    .R(_01944_),
    .S(1'h1)
  );
  DFFSR _10016_ (
    .CLK(dco_clk),
    .D(_02176_),
    .Q( execution_unit_0.register_file_0.r13_6_ ),
    .R(_01945_),
    .S(1'h1)
  );
  DFFSR _10017_ (
    .CLK(dco_clk),
    .D(_02177_),
    .Q( execution_unit_0.register_file_0.r13_7_ ),
    .R(_01946_),
    .S(1'h1)
  );
  DFFSR _10018_ (
    .CLK(dco_clk),
    .D(_02178_),
    .Q( execution_unit_0.register_file_0.r13_8_ ),
    .R(_01947_),
    .S(1'h1)
  );
  DFFSR _10019_ (
    .CLK(dco_clk),
    .D(_02179_),
    .Q( execution_unit_0.register_file_0.r13_9_ ),
    .R(_01948_),
    .S(1'h1)
  );
  DFFSR _10020_ (
    .CLK(dco_clk),
    .D(_02180_),
    .Q( execution_unit_0.register_file_0.r13_10_ ),
    .R(_01949_),
    .S(1'h1)
  );
  DFFSR _10021_ (
    .CLK(dco_clk),
    .D(_02181_),
    .Q( execution_unit_0.register_file_0.r13_11_ ),
    .R(_01950_),
    .S(1'h1)
  );
  DFFSR _10022_ (
    .CLK(dco_clk),
    .D(_02182_),
    .Q( execution_unit_0.register_file_0.r13_12_ ),
    .R(_01951_),
    .S(1'h1)
  );
  DFFSR _10023_ (
    .CLK(dco_clk),
    .D(_02183_),
    .Q( execution_unit_0.register_file_0.r13_13_ ),
    .R(_01952_),
    .S(1'h1)
  );
  DFFSR _10024_ (
    .CLK(dco_clk),
    .D(_02184_),
    .Q( execution_unit_0.register_file_0.r13_14_ ),
    .R(_01953_),
    .S(1'h1)
  );
  DFFSR _10025_ (
    .CLK(dco_clk),
    .D(_02185_),
    .Q( execution_unit_0.register_file_0.r13_15_ ),
    .R(_01954_),
    .S(1'h1)
  );
  DFFSR _10026_ (
    .CLK(dco_clk),
    .D(_02186_),
    .Q( execution_unit_0.register_file_0.r12_0_ ),
    .R(_01955_),
    .S(1'h1)
  );
  DFFSR _10027_ (
    .CLK(dco_clk),
    .D(_02187_),
    .Q( execution_unit_0.register_file_0.r12_1_ ),
    .R(_01956_),
    .S(1'h1)
  );
  DFFSR _10028_ (
    .CLK(dco_clk),
    .D(_02188_),
    .Q( execution_unit_0.register_file_0.r12_2_ ),
    .R(_01957_),
    .S(1'h1)
  );
  DFFSR _10029_ (
    .CLK(dco_clk),
    .D(_02189_),
    .Q( execution_unit_0.register_file_0.r12_3_ ),
    .R(_01958_),
    .S(1'h1)
  );
  DFFSR _10030_ (
    .CLK(dco_clk),
    .D(_02190_),
    .Q( execution_unit_0.register_file_0.r12_4_ ),
    .R(_01959_),
    .S(1'h1)
  );
  DFFSR _10031_ (
    .CLK(dco_clk),
    .D(_02191_),
    .Q( execution_unit_0.register_file_0.r12_5_ ),
    .R(_01960_),
    .S(1'h1)
  );
  DFFSR _10032_ (
    .CLK(dco_clk),
    .D(_02192_),
    .Q( execution_unit_0.register_file_0.r12_6_ ),
    .R(_01961_),
    .S(1'h1)
  );
  DFFSR _10033_ (
    .CLK(dco_clk),
    .D(_02193_),
    .Q( execution_unit_0.register_file_0.r12_7_ ),
    .R(_01962_),
    .S(1'h1)
  );
  DFFSR _10034_ (
    .CLK(dco_clk),
    .D(_02194_),
    .Q( execution_unit_0.register_file_0.r12_8_ ),
    .R(_01963_),
    .S(1'h1)
  );
  DFFSR _10035_ (
    .CLK(dco_clk),
    .D(_02195_),
    .Q( execution_unit_0.register_file_0.r12_9_ ),
    .R(_01964_),
    .S(1'h1)
  );
  DFFSR _10036_ (
    .CLK(dco_clk),
    .D(_02196_),
    .Q( execution_unit_0.register_file_0.r12_10_ ),
    .R(_01965_),
    .S(1'h1)
  );
  DFFSR _10037_ (
    .CLK(dco_clk),
    .D(_02197_),
    .Q( execution_unit_0.register_file_0.r12_11_ ),
    .R(_01966_),
    .S(1'h1)
  );
  DFFSR _10038_ (
    .CLK(dco_clk),
    .D(_02198_),
    .Q( execution_unit_0.register_file_0.r12_12_ ),
    .R(_01967_),
    .S(1'h1)
  );
  DFFSR _10039_ (
    .CLK(dco_clk),
    .D(_02199_),
    .Q( execution_unit_0.register_file_0.r12_13_ ),
    .R(_01968_),
    .S(1'h1)
  );
  DFFSR _10040_ (
    .CLK(dco_clk),
    .D(_02200_),
    .Q( execution_unit_0.register_file_0.r12_14_ ),
    .R(_01969_),
    .S(1'h1)
  );
  DFFSR _10041_ (
    .CLK(dco_clk),
    .D(_02201_),
    .Q( execution_unit_0.register_file_0.r12_15_ ),
    .R(_01970_),
    .S(1'h1)
  );
  DFFSR _10042_ (
    .CLK(dco_clk),
    .D(_02202_),
    .Q( execution_unit_0.register_file_0.r11_0_ ),
    .R(_01971_),
    .S(1'h1)
  );
  DFFSR _10043_ (
    .CLK(dco_clk),
    .D(_02203_),
    .Q( execution_unit_0.register_file_0.r11_1_ ),
    .R(_01972_),
    .S(1'h1)
  );
  DFFSR _10044_ (
    .CLK(dco_clk),
    .D(_02204_),
    .Q( execution_unit_0.register_file_0.r11_2_ ),
    .R(_01973_),
    .S(1'h1)
  );
  DFFSR _10045_ (
    .CLK(dco_clk),
    .D(_02205_),
    .Q( execution_unit_0.register_file_0.r11_3_ ),
    .R(_01974_),
    .S(1'h1)
  );
  DFFSR _10046_ (
    .CLK(dco_clk),
    .D(_02206_),
    .Q( execution_unit_0.register_file_0.r11_4_ ),
    .R(_01975_),
    .S(1'h1)
  );
  DFFSR _10047_ (
    .CLK(dco_clk),
    .D(_02207_),
    .Q( execution_unit_0.register_file_0.r11_5_ ),
    .R(_01976_),
    .S(1'h1)
  );
  DFFSR _10048_ (
    .CLK(dco_clk),
    .D(_02208_),
    .Q( execution_unit_0.register_file_0.r11_6_ ),
    .R(_01977_),
    .S(1'h1)
  );
  DFFSR _10049_ (
    .CLK(dco_clk),
    .D(_02209_),
    .Q( execution_unit_0.register_file_0.r11_7_ ),
    .R(_01978_),
    .S(1'h1)
  );
  DFFSR _10050_ (
    .CLK(dco_clk),
    .D(_02210_),
    .Q( execution_unit_0.register_file_0.r11_8_ ),
    .R(_01979_),
    .S(1'h1)
  );
  DFFSR _10051_ (
    .CLK(dco_clk),
    .D(_02211_),
    .Q( execution_unit_0.register_file_0.r11_9_ ),
    .R(_01980_),
    .S(1'h1)
  );
  DFFSR _10052_ (
    .CLK(dco_clk),
    .D(_02212_),
    .Q( execution_unit_0.register_file_0.r11_10_ ),
    .R(_01981_),
    .S(1'h1)
  );
  DFFSR _10053_ (
    .CLK(dco_clk),
    .D(_02213_),
    .Q( execution_unit_0.register_file_0.r11_11_ ),
    .R(_01982_),
    .S(1'h1)
  );
  DFFSR _10054_ (
    .CLK(dco_clk),
    .D(_02214_),
    .Q( execution_unit_0.register_file_0.r11_12_ ),
    .R(_01983_),
    .S(1'h1)
  );
  DFFSR _10055_ (
    .CLK(dco_clk),
    .D(_02215_),
    .Q( execution_unit_0.register_file_0.r11_13_ ),
    .R(_01984_),
    .S(1'h1)
  );
  DFFSR _10056_ (
    .CLK(dco_clk),
    .D(_02216_),
    .Q( execution_unit_0.register_file_0.r11_14_ ),
    .R(_01985_),
    .S(1'h1)
  );
  DFFSR _10057_ (
    .CLK(dco_clk),
    .D(_02217_),
    .Q( execution_unit_0.register_file_0.r11_15_ ),
    .R(_01986_),
    .S(1'h1)
  );
  DFFSR _10058_ (
    .CLK(dco_clk),
    .D(_02218_),
    .Q( execution_unit_0.register_file_0.r10_0_ ),
    .R(_01987_),
    .S(1'h1)
  );
  DFFSR _10059_ (
    .CLK(dco_clk),
    .D(_02219_),
    .Q( execution_unit_0.register_file_0.r10_1_ ),
    .R(_01988_),
    .S(1'h1)
  );
  DFFSR _10060_ (
    .CLK(dco_clk),
    .D(_02220_),
    .Q( execution_unit_0.register_file_0.r10_2_ ),
    .R(_01989_),
    .S(1'h1)
  );
  DFFSR _10061_ (
    .CLK(dco_clk),
    .D(_02221_),
    .Q( execution_unit_0.register_file_0.r10_3_ ),
    .R(_01990_),
    .S(1'h1)
  );
  DFFSR _10062_ (
    .CLK(dco_clk),
    .D(_02222_),
    .Q( execution_unit_0.register_file_0.r10_4_ ),
    .R(_01991_),
    .S(1'h1)
  );
  DFFSR _10063_ (
    .CLK(dco_clk),
    .D(_02223_),
    .Q( execution_unit_0.register_file_0.r10_5_ ),
    .R(_01992_),
    .S(1'h1)
  );
  DFFSR _10064_ (
    .CLK(dco_clk),
    .D(_02224_),
    .Q( execution_unit_0.register_file_0.r10_6_ ),
    .R(_01993_),
    .S(1'h1)
  );
  DFFSR _10065_ (
    .CLK(dco_clk),
    .D(_02225_),
    .Q( execution_unit_0.register_file_0.r10_7_ ),
    .R(_01994_),
    .S(1'h1)
  );
  DFFSR _10066_ (
    .CLK(dco_clk),
    .D(_02226_),
    .Q( execution_unit_0.register_file_0.r10_8_ ),
    .R(_01995_),
    .S(1'h1)
  );
  DFFSR _10067_ (
    .CLK(dco_clk),
    .D(_02227_),
    .Q( execution_unit_0.register_file_0.r10_9_ ),
    .R(_01996_),
    .S(1'h1)
  );
  DFFSR _10068_ (
    .CLK(dco_clk),
    .D(_02228_),
    .Q( execution_unit_0.register_file_0.r10_10_ ),
    .R(_01997_),
    .S(1'h1)
  );
  DFFSR _10069_ (
    .CLK(dco_clk),
    .D(_02229_),
    .Q( execution_unit_0.register_file_0.r10_11_ ),
    .R(_01998_),
    .S(1'h1)
  );
  DFFSR _10070_ (
    .CLK(dco_clk),
    .D(_02230_),
    .Q( execution_unit_0.register_file_0.r10_12_ ),
    .R(_01999_),
    .S(1'h1)
  );
  DFFSR _10071_ (
    .CLK(dco_clk),
    .D(_02231_),
    .Q( execution_unit_0.register_file_0.r10_13_ ),
    .R(_02000_),
    .S(1'h1)
  );
  DFFSR _10072_ (
    .CLK(dco_clk),
    .D(_02232_),
    .Q( execution_unit_0.register_file_0.r10_14_ ),
    .R(_02001_),
    .S(1'h1)
  );
  DFFSR _10073_ (
    .CLK(dco_clk),
    .D(_02233_),
    .Q( execution_unit_0.register_file_0.r10_15_ ),
    .R(_02002_),
    .S(1'h1)
  );
  DFFSR _10074_ (
    .CLK(dco_clk),
    .D(_02234_),
    .Q( execution_unit_0.register_file_0.r9_0_ ),
    .R(_02003_),
    .S(1'h1)
  );
  DFFSR _10075_ (
    .CLK(dco_clk),
    .D(_02235_),
    .Q( execution_unit_0.register_file_0.r9_1_ ),
    .R(_02004_),
    .S(1'h1)
  );
  DFFSR _10076_ (
    .CLK(dco_clk),
    .D(_02236_),
    .Q( execution_unit_0.register_file_0.r9_2_ ),
    .R(_02005_),
    .S(1'h1)
  );
  DFFSR _10077_ (
    .CLK(dco_clk),
    .D(_02237_),
    .Q( execution_unit_0.register_file_0.r9_3_ ),
    .R(_02006_),
    .S(1'h1)
  );
  DFFSR _10078_ (
    .CLK(dco_clk),
    .D(_02238_),
    .Q( execution_unit_0.register_file_0.r9_4_ ),
    .R(_02007_),
    .S(1'h1)
  );
  DFFSR _10079_ (
    .CLK(dco_clk),
    .D(_02239_),
    .Q( execution_unit_0.register_file_0.r9_5_ ),
    .R(_02008_),
    .S(1'h1)
  );
  DFFSR _10080_ (
    .CLK(dco_clk),
    .D(_02240_),
    .Q( execution_unit_0.register_file_0.r9_6_ ),
    .R(_02009_),
    .S(1'h1)
  );
  DFFSR _10081_ (
    .CLK(dco_clk),
    .D(_02241_),
    .Q( execution_unit_0.register_file_0.r9_7_ ),
    .R(_02010_),
    .S(1'h1)
  );
  DFFSR _10082_ (
    .CLK(dco_clk),
    .D(_02242_),
    .Q( execution_unit_0.register_file_0.r9_8_ ),
    .R(_02011_),
    .S(1'h1)
  );
  DFFSR _10083_ (
    .CLK(dco_clk),
    .D(_02243_),
    .Q( execution_unit_0.register_file_0.r9_9_ ),
    .R(_02012_),
    .S(1'h1)
  );
  DFFSR _10084_ (
    .CLK(dco_clk),
    .D(_02244_),
    .Q( execution_unit_0.register_file_0.r9_10_ ),
    .R(_02013_),
    .S(1'h1)
  );
  DFFSR _10085_ (
    .CLK(dco_clk),
    .D(_02245_),
    .Q( execution_unit_0.register_file_0.r9_11_ ),
    .R(_02014_),
    .S(1'h1)
  );
  DFFSR _10086_ (
    .CLK(dco_clk),
    .D(_02246_),
    .Q( execution_unit_0.register_file_0.r9_12_ ),
    .R(_02015_),
    .S(1'h1)
  );
  DFFSR _10087_ (
    .CLK(dco_clk),
    .D(_02247_),
    .Q( execution_unit_0.register_file_0.r9_13_ ),
    .R(_02016_),
    .S(1'h1)
  );
  DFFSR _10088_ (
    .CLK(dco_clk),
    .D(_02248_),
    .Q( execution_unit_0.register_file_0.r9_14_ ),
    .R(_02017_),
    .S(1'h1)
  );
  DFFSR _10089_ (
    .CLK(dco_clk),
    .D(_02249_),
    .Q( execution_unit_0.register_file_0.r9_15_ ),
    .R(_02018_),
    .S(1'h1)
  );
  DFFSR _10090_ (
    .CLK(dco_clk),
    .D(_02250_),
    .Q( execution_unit_0.register_file_0.r8_0_ ),
    .R(_02019_),
    .S(1'h1)
  );
  DFFSR _10091_ (
    .CLK(dco_clk),
    .D(_02251_),
    .Q( execution_unit_0.register_file_0.r8_1_ ),
    .R(_02020_),
    .S(1'h1)
  );
  DFFSR _10092_ (
    .CLK(dco_clk),
    .D(_02252_),
    .Q( execution_unit_0.register_file_0.r8_2_ ),
    .R(_02021_),
    .S(1'h1)
  );
  DFFSR _10093_ (
    .CLK(dco_clk),
    .D(_02253_),
    .Q( execution_unit_0.register_file_0.r8_3_ ),
    .R(_02022_),
    .S(1'h1)
  );
  DFFSR _10094_ (
    .CLK(dco_clk),
    .D(_02254_),
    .Q( execution_unit_0.register_file_0.r8_4_ ),
    .R(_02023_),
    .S(1'h1)
  );
  DFFSR _10095_ (
    .CLK(dco_clk),
    .D(_02255_),
    .Q( execution_unit_0.register_file_0.r8_5_ ),
    .R(_02024_),
    .S(1'h1)
  );
  DFFSR _10096_ (
    .CLK(dco_clk),
    .D(_02256_),
    .Q( execution_unit_0.register_file_0.r8_6_ ),
    .R(_02025_),
    .S(1'h1)
  );
  DFFSR _10097_ (
    .CLK(dco_clk),
    .D(_02257_),
    .Q( execution_unit_0.register_file_0.r8_7_ ),
    .R(_02026_),
    .S(1'h1)
  );
  DFFSR _10098_ (
    .CLK(dco_clk),
    .D(_02258_),
    .Q( execution_unit_0.register_file_0.r8_8_ ),
    .R(_02027_),
    .S(1'h1)
  );
  DFFSR _10099_ (
    .CLK(dco_clk),
    .D(_02259_),
    .Q( execution_unit_0.register_file_0.r8_9_ ),
    .R(_02028_),
    .S(1'h1)
  );
  DFFSR _10100_ (
    .CLK(dco_clk),
    .D(_02260_),
    .Q( execution_unit_0.register_file_0.r8_10_ ),
    .R(_02029_),
    .S(1'h1)
  );
  DFFSR _10101_ (
    .CLK(dco_clk),
    .D(_02261_),
    .Q( execution_unit_0.register_file_0.r8_11_ ),
    .R(_02030_),
    .S(1'h1)
  );
  DFFSR _10102_ (
    .CLK(dco_clk),
    .D(_02262_),
    .Q( execution_unit_0.register_file_0.r8_12_ ),
    .R(_02031_),
    .S(1'h1)
  );
  DFFSR _10103_ (
    .CLK(dco_clk),
    .D(_02263_),
    .Q( execution_unit_0.register_file_0.r8_13_ ),
    .R(_02032_),
    .S(1'h1)
  );
  DFFSR _10104_ (
    .CLK(dco_clk),
    .D(_02264_),
    .Q( execution_unit_0.register_file_0.r8_14_ ),
    .R(_02033_),
    .S(1'h1)
  );
  DFFSR _10105_ (
    .CLK(dco_clk),
    .D(_02265_),
    .Q( execution_unit_0.register_file_0.r8_15_ ),
    .R(_02034_),
    .S(1'h1)
  );
  DFFSR _10106_ (
    .CLK(dco_clk),
    .D(_02266_),
    .Q( execution_unit_0.register_file_0.r7_0_ ),
    .R(_02035_),
    .S(1'h1)
  );
  DFFSR _10107_ (
    .CLK(dco_clk),
    .D(_02267_),
    .Q( execution_unit_0.register_file_0.r7_1_ ),
    .R(_02036_),
    .S(1'h1)
  );
  DFFSR _10108_ (
    .CLK(dco_clk),
    .D(_02268_),
    .Q( execution_unit_0.register_file_0.r7_2_ ),
    .R(_02037_),
    .S(1'h1)
  );
  DFFSR _10109_ (
    .CLK(dco_clk),
    .D(_02269_),
    .Q( execution_unit_0.register_file_0.r7_3_ ),
    .R(_02038_),
    .S(1'h1)
  );
  DFFSR _10110_ (
    .CLK(dco_clk),
    .D(_02270_),
    .Q( execution_unit_0.register_file_0.r7_4_ ),
    .R(_02039_),
    .S(1'h1)
  );
  DFFSR _10111_ (
    .CLK(dco_clk),
    .D(_02271_),
    .Q( execution_unit_0.register_file_0.r7_5_ ),
    .R(_02040_),
    .S(1'h1)
  );
  DFFSR _10112_ (
    .CLK(dco_clk),
    .D(_02272_),
    .Q( execution_unit_0.register_file_0.r7_6_ ),
    .R(_02041_),
    .S(1'h1)
  );
  DFFSR _10113_ (
    .CLK(dco_clk),
    .D(_02273_),
    .Q( execution_unit_0.register_file_0.r7_7_ ),
    .R(_02042_),
    .S(1'h1)
  );
  DFFSR _10114_ (
    .CLK(dco_clk),
    .D(_02274_),
    .Q( execution_unit_0.register_file_0.r7_8_ ),
    .R(_02043_),
    .S(1'h1)
  );
  DFFSR _10115_ (
    .CLK(dco_clk),
    .D(_02275_),
    .Q( execution_unit_0.register_file_0.r7_9_ ),
    .R(_02044_),
    .S(1'h1)
  );
  DFFSR _10116_ (
    .CLK(dco_clk),
    .D(_02276_),
    .Q( execution_unit_0.register_file_0.r7_10_ ),
    .R(_02045_),
    .S(1'h1)
  );
  DFFSR _10117_ (
    .CLK(dco_clk),
    .D(_02277_),
    .Q( execution_unit_0.register_file_0.r7_11_ ),
    .R(_02046_),
    .S(1'h1)
  );
  DFFSR _10118_ (
    .CLK(dco_clk),
    .D(_02278_),
    .Q( execution_unit_0.register_file_0.r7_12_ ),
    .R(_02047_),
    .S(1'h1)
  );
  DFFSR _10119_ (
    .CLK(dco_clk),
    .D(_02279_),
    .Q( execution_unit_0.register_file_0.r7_13_ ),
    .R(_02048_),
    .S(1'h1)
  );
  DFFSR _10120_ (
    .CLK(dco_clk),
    .D(_02280_),
    .Q( execution_unit_0.register_file_0.r7_14_ ),
    .R(_02049_),
    .S(1'h1)
  );
  DFFSR _10121_ (
    .CLK(dco_clk),
    .D(_02281_),
    .Q( execution_unit_0.register_file_0.r7_15_ ),
    .R(_02050_),
    .S(1'h1)
  );
  DFFSR _10122_ (
    .CLK(dco_clk),
    .D(_02282_),
    .Q( execution_unit_0.register_file_0.r6_0_ ),
    .R(_02051_),
    .S(1'h1)
  );
  DFFSR _10123_ (
    .CLK(dco_clk),
    .D(_02283_),
    .Q( execution_unit_0.register_file_0.r6_1_ ),
    .R(_02052_),
    .S(1'h1)
  );
  DFFSR _10124_ (
    .CLK(dco_clk),
    .D(_02284_),
    .Q( execution_unit_0.register_file_0.r6_2_ ),
    .R(_02053_),
    .S(1'h1)
  );
  DFFSR _10125_ (
    .CLK(dco_clk),
    .D(_02285_),
    .Q( execution_unit_0.register_file_0.r6_3_ ),
    .R(_02054_),
    .S(1'h1)
  );
  DFFSR _10126_ (
    .CLK(dco_clk),
    .D(_02286_),
    .Q( execution_unit_0.register_file_0.r6_4_ ),
    .R(_02055_),
    .S(1'h1)
  );
  DFFSR _10127_ (
    .CLK(dco_clk),
    .D(_02287_),
    .Q( execution_unit_0.register_file_0.r6_5_ ),
    .R(_02056_),
    .S(1'h1)
  );
  DFFSR _10128_ (
    .CLK(dco_clk),
    .D(_02288_),
    .Q( execution_unit_0.register_file_0.r6_6_ ),
    .R(_02057_),
    .S(1'h1)
  );
  DFFSR _10129_ (
    .CLK(dco_clk),
    .D(_02289_),
    .Q( execution_unit_0.register_file_0.r6_7_ ),
    .R(_02058_),
    .S(1'h1)
  );
  DFFSR _10130_ (
    .CLK(dco_clk),
    .D(_02290_),
    .Q( execution_unit_0.register_file_0.r6_8_ ),
    .R(_02059_),
    .S(1'h1)
  );
  DFFSR _10131_ (
    .CLK(dco_clk),
    .D(_02291_),
    .Q( execution_unit_0.register_file_0.r6_9_ ),
    .R(_02060_),
    .S(1'h1)
  );
  DFFSR _10132_ (
    .CLK(dco_clk),
    .D(_02292_),
    .Q( execution_unit_0.register_file_0.r6_10_ ),
    .R(_02061_),
    .S(1'h1)
  );
  DFFSR _10133_ (
    .CLK(dco_clk),
    .D(_02293_),
    .Q( execution_unit_0.register_file_0.r6_11_ ),
    .R(_02062_),
    .S(1'h1)
  );
  DFFSR _10134_ (
    .CLK(dco_clk),
    .D(_02294_),
    .Q( execution_unit_0.register_file_0.r6_12_ ),
    .R(_02063_),
    .S(1'h1)
  );
  DFFSR _10135_ (
    .CLK(dco_clk),
    .D(_02295_),
    .Q( execution_unit_0.register_file_0.r6_13_ ),
    .R(_02064_),
    .S(1'h1)
  );
  DFFSR _10136_ (
    .CLK(dco_clk),
    .D(_02296_),
    .Q( execution_unit_0.register_file_0.r6_14_ ),
    .R(_02065_),
    .S(1'h1)
  );
  DFFSR _10137_ (
    .CLK(dco_clk),
    .D(_02297_),
    .Q( execution_unit_0.register_file_0.r6_15_ ),
    .R(_02066_),
    .S(1'h1)
  );
  DFFSR _10138_ (
    .CLK(dco_clk),
    .D(_02298_),
    .Q( execution_unit_0.register_file_0.r5_0_ ),
    .R(_02067_),
    .S(1'h1)
  );
  DFFSR _10139_ (
    .CLK(dco_clk),
    .D(_02299_),
    .Q( execution_unit_0.register_file_0.r5_1_ ),
    .R(_02068_),
    .S(1'h1)
  );
  DFFSR _10140_ (
    .CLK(dco_clk),
    .D(_02300_),
    .Q( execution_unit_0.register_file_0.r5_2_ ),
    .R(_02069_),
    .S(1'h1)
  );
  DFFSR _10141_ (
    .CLK(dco_clk),
    .D(_02301_),
    .Q( execution_unit_0.register_file_0.r5_3_ ),
    .R(_02070_),
    .S(1'h1)
  );
  DFFSR _10142_ (
    .CLK(dco_clk),
    .D(_02302_),
    .Q( execution_unit_0.register_file_0.r5_4_ ),
    .R(_02071_),
    .S(1'h1)
  );
  DFFSR _10143_ (
    .CLK(dco_clk),
    .D(_02303_),
    .Q( execution_unit_0.register_file_0.r5_5_ ),
    .R(_02072_),
    .S(1'h1)
  );
  DFFSR _10144_ (
    .CLK(dco_clk),
    .D(_02304_),
    .Q( execution_unit_0.register_file_0.r5_6_ ),
    .R(_02073_),
    .S(1'h1)
  );
  DFFSR _10145_ (
    .CLK(dco_clk),
    .D(_02305_),
    .Q( execution_unit_0.register_file_0.r5_7_ ),
    .R(_02074_),
    .S(1'h1)
  );
  DFFSR _10146_ (
    .CLK(dco_clk),
    .D(_02306_),
    .Q( execution_unit_0.register_file_0.r5_8_ ),
    .R(_02075_),
    .S(1'h1)
  );
  DFFSR _10147_ (
    .CLK(dco_clk),
    .D(_02307_),
    .Q( execution_unit_0.register_file_0.r5_9_ ),
    .R(_02076_),
    .S(1'h1)
  );
  DFFSR _10148_ (
    .CLK(dco_clk),
    .D(_02308_),
    .Q( execution_unit_0.register_file_0.r5_10_ ),
    .R(_02077_),
    .S(1'h1)
  );
  DFFSR _10149_ (
    .CLK(dco_clk),
    .D(_02309_),
    .Q( execution_unit_0.register_file_0.r5_11_ ),
    .R(_02078_),
    .S(1'h1)
  );
  DFFSR _10150_ (
    .CLK(dco_clk),
    .D(_02310_),
    .Q( execution_unit_0.register_file_0.r5_12_ ),
    .R(_02079_),
    .S(1'h1)
  );
  DFFSR _10151_ (
    .CLK(dco_clk),
    .D(_02311_),
    .Q( execution_unit_0.register_file_0.r5_13_ ),
    .R(_02080_),
    .S(1'h1)
  );
  DFFSR _10152_ (
    .CLK(dco_clk),
    .D(_02312_),
    .Q( execution_unit_0.register_file_0.r5_14_ ),
    .R(_02081_),
    .S(1'h1)
  );
  DFFSR _10153_ (
    .CLK(dco_clk),
    .D(_02313_),
    .Q( execution_unit_0.register_file_0.r5_15_ ),
    .R(_02082_),
    .S(1'h1)
  );
  DFFSR _10154_ (
    .CLK(dco_clk),
    .D(_02314_),
    .Q( execution_unit_0.register_file_0.r4_0_ ),
    .R(_02083_),
    .S(1'h1)
  );
  DFFSR _10155_ (
    .CLK(dco_clk),
    .D(_02315_),
    .Q( execution_unit_0.register_file_0.r4_1_ ),
    .R(_02084_),
    .S(1'h1)
  );
  DFFSR _10156_ (
    .CLK(dco_clk),
    .D(_02316_),
    .Q( execution_unit_0.register_file_0.r4_2_ ),
    .R(_02085_),
    .S(1'h1)
  );
  DFFSR _10157_ (
    .CLK(dco_clk),
    .D(_02317_),
    .Q( execution_unit_0.register_file_0.r4_3_ ),
    .R(_02086_),
    .S(1'h1)
  );
  DFFSR _10158_ (
    .CLK(dco_clk),
    .D(_02318_),
    .Q( execution_unit_0.register_file_0.r4_4_ ),
    .R(_02087_),
    .S(1'h1)
  );
  DFFSR _10159_ (
    .CLK(dco_clk),
    .D(_02319_),
    .Q( execution_unit_0.register_file_0.r4_5_ ),
    .R(_02088_),
    .S(1'h1)
  );
  DFFSR _10160_ (
    .CLK(dco_clk),
    .D(_02320_),
    .Q( execution_unit_0.register_file_0.r4_6_ ),
    .R(_02089_),
    .S(1'h1)
  );
  DFFSR _10161_ (
    .CLK(dco_clk),
    .D(_02321_),
    .Q( execution_unit_0.register_file_0.r4_7_ ),
    .R(_02090_),
    .S(1'h1)
  );
  DFFSR _10162_ (
    .CLK(dco_clk),
    .D(_02322_),
    .Q( execution_unit_0.register_file_0.r4_8_ ),
    .R(_02091_),
    .S(1'h1)
  );
  DFFSR _10163_ (
    .CLK(dco_clk),
    .D(_02323_),
    .Q( execution_unit_0.register_file_0.r4_9_ ),
    .R(_02092_),
    .S(1'h1)
  );
  DFFSR _10164_ (
    .CLK(dco_clk),
    .D(_02324_),
    .Q( execution_unit_0.register_file_0.r4_10_ ),
    .R(_02093_),
    .S(1'h1)
  );
  DFFSR _10165_ (
    .CLK(dco_clk),
    .D(_02325_),
    .Q( execution_unit_0.register_file_0.r4_11_ ),
    .R(_02094_),
    .S(1'h1)
  );
  DFFSR _10166_ (
    .CLK(dco_clk),
    .D(_02326_),
    .Q( execution_unit_0.register_file_0.r4_12_ ),
    .R(_02095_),
    .S(1'h1)
  );
  DFFSR _10167_ (
    .CLK(dco_clk),
    .D(_02327_),
    .Q( execution_unit_0.register_file_0.r4_13_ ),
    .R(_02096_),
    .S(1'h1)
  );
  DFFSR _10168_ (
    .CLK(dco_clk),
    .D(_02328_),
    .Q( execution_unit_0.register_file_0.r4_14_ ),
    .R(_02097_),
    .S(1'h1)
  );
  DFFSR _10169_ (
    .CLK(dco_clk),
    .D(_02329_),
    .Q( execution_unit_0.register_file_0.r4_15_ ),
    .R(_02098_),
    .S(1'h1)
  );
  DFFSR _10170_ (
    .CLK(dco_clk),
    .D(_02330_),
    .Q( execution_unit_0.register_file_0.r3_0_ ),
    .R(_02099_),
    .S(1'h1)
  );
  DFFSR _10171_ (
    .CLK(dco_clk),
    .D(_02331_),
    .Q( execution_unit_0.register_file_0.r3_1_ ),
    .R(_02100_),
    .S(1'h1)
  );
  DFFSR _10172_ (
    .CLK(dco_clk),
    .D(_02332_),
    .Q( execution_unit_0.register_file_0.r3_2_ ),
    .R(_02101_),
    .S(1'h1)
  );
  DFFSR _10173_ (
    .CLK(dco_clk),
    .D(_02333_),
    .Q( execution_unit_0.register_file_0.r3_3_ ),
    .R(_02102_),
    .S(1'h1)
  );
  DFFSR _10174_ (
    .CLK(dco_clk),
    .D(_02334_),
    .Q( execution_unit_0.register_file_0.r3_4_ ),
    .R(_02103_),
    .S(1'h1)
  );
  DFFSR _10175_ (
    .CLK(dco_clk),
    .D(_02335_),
    .Q( execution_unit_0.register_file_0.r3_5_ ),
    .R(_02104_),
    .S(1'h1)
  );
  DFFSR _10176_ (
    .CLK(dco_clk),
    .D(_02336_),
    .Q( execution_unit_0.register_file_0.r3_6_ ),
    .R(_02105_),
    .S(1'h1)
  );
  DFFSR _10177_ (
    .CLK(dco_clk),
    .D(_02337_),
    .Q( execution_unit_0.register_file_0.r3_7_ ),
    .R(_02106_),
    .S(1'h1)
  );
  DFFSR _10178_ (
    .CLK(dco_clk),
    .D(_02338_),
    .Q( execution_unit_0.register_file_0.r3_8_ ),
    .R(_02107_),
    .S(1'h1)
  );
  DFFSR _10179_ (
    .CLK(dco_clk),
    .D(_02339_),
    .Q( execution_unit_0.register_file_0.r3_9_ ),
    .R(_02108_),
    .S(1'h1)
  );
  DFFSR _10180_ (
    .CLK(dco_clk),
    .D(_02340_),
    .Q( execution_unit_0.register_file_0.r3_10_ ),
    .R(_02109_),
    .S(1'h1)
  );
  DFFSR _10181_ (
    .CLK(dco_clk),
    .D(_02341_),
    .Q( execution_unit_0.register_file_0.r3_11_ ),
    .R(_02110_),
    .S(1'h1)
  );
  DFFSR _10182_ (
    .CLK(dco_clk),
    .D(_02342_),
    .Q( execution_unit_0.register_file_0.r3_12_ ),
    .R(_02111_),
    .S(1'h1)
  );
  DFFSR _10183_ (
    .CLK(dco_clk),
    .D(_02343_),
    .Q( execution_unit_0.register_file_0.r3_13_ ),
    .R(_02112_),
    .S(1'h1)
  );
  DFFSR _10184_ (
    .CLK(dco_clk),
    .D(_02344_),
    .Q( execution_unit_0.register_file_0.r3_14_ ),
    .R(_02113_),
    .S(1'h1)
  );
  DFFSR _10185_ (
    .CLK(dco_clk),
    .D(_02345_),
    .Q( execution_unit_0.register_file_0.r3_15_ ),
    .R(_02114_),
    .S(1'h1)
  );
  DFFSR _10186_ (
    .CLK(dco_clk),
    .D(_02346_),
    .Q( execution_unit_0.alu_0.status_0_ ),
    .R(_02115_),
    .S(1'h1)
  );
  DFFSR _10187_ (
    .CLK(dco_clk),
    .D(_01900_),
    .Q( execution_unit_0.register_file_0.r2_4_ ),
    .R(_02116_),
    .S(1'h1)
  );
  DFFSR _10188_ (
    .CLK(dco_clk),
    .D(_02347_),
    .Q( execution_unit_0.register_file_0.r1_1_ ),
    .R(_02117_),
    .S(1'h1)
  );
  DFFSR _10189_ (
    .CLK(dco_clk),
    .D(_02348_),
    .Q( execution_unit_0.register_file_0.r1_2_ ),
    .R(_02118_),
    .S(1'h1)
  );
  DFFSR _10190_ (
    .CLK(dco_clk),
    .D(_02349_),
    .Q( execution_unit_0.register_file_0.r1_3_ ),
    .R(_02119_),
    .S(1'h1)
  );
  DFFSR _10191_ (
    .CLK(dco_clk),
    .D(_02350_),
    .Q( execution_unit_0.register_file_0.r1_4_ ),
    .R(_02120_),
    .S(1'h1)
  );
  DFFSR _10192_ (
    .CLK(dco_clk),
    .D(_02351_),
    .Q( execution_unit_0.register_file_0.r1_5_ ),
    .R(_02121_),
    .S(1'h1)
  );
  DFFSR _10193_ (
    .CLK(dco_clk),
    .D(_02352_),
    .Q( execution_unit_0.register_file_0.r1_6_ ),
    .R(_02122_),
    .S(1'h1)
  );
  DFFSR _10194_ (
    .CLK(dco_clk),
    .D(_02353_),
    .Q( execution_unit_0.register_file_0.r1_7_ ),
    .R(_02123_),
    .S(1'h1)
  );
  DFFSR _10195_ (
    .CLK(dco_clk),
    .D(_02354_),
    .Q( execution_unit_0.register_file_0.r1_8_ ),
    .R(_02124_),
    .S(1'h1)
  );
  DFFSR _10196_ (
    .CLK(dco_clk),
    .D(_02355_),
    .Q( execution_unit_0.register_file_0.r1_9_ ),
    .R(_02125_),
    .S(1'h1)
  );
  DFFSR _10197_ (
    .CLK(dco_clk),
    .D(_02356_),
    .Q( execution_unit_0.register_file_0.r1_10_ ),
    .R(_02126_),
    .S(1'h1)
  );
  DFFSR _10198_ (
    .CLK(dco_clk),
    .D(_02357_),
    .Q( execution_unit_0.register_file_0.r1_11_ ),
    .R(_02127_),
    .S(1'h1)
  );
  DFFSR _10199_ (
    .CLK(dco_clk),
    .D(_02358_),
    .Q( execution_unit_0.register_file_0.r1_12_ ),
    .R(_02128_),
    .S(1'h1)
  );
  DFFSR _10200_ (
    .CLK(dco_clk),
    .D(_02359_),
    .Q( execution_unit_0.register_file_0.r1_13_ ),
    .R(_02129_),
    .S(1'h1)
  );
  DFFSR _10201_ (
    .CLK(dco_clk),
    .D(_02360_),
    .Q( execution_unit_0.register_file_0.r1_14_ ),
    .R(_02130_),
    .S(1'h1)
  );
  DFFSR _10202_ (
    .CLK(dco_clk),
    .D(_02361_),
    .Q( execution_unit_0.register_file_0.r1_15_ ),
    .R(_02131_),
    .S(1'h1)
  );
  INVX1 _10203_ (
    .A( frontend_0.irq_addr_3_ ),
    .Y(_03743_)
  );
  INVX1 _10204_ (
    .A( frontend_0.irq_addr_2_ ),
    .Y(_03744_)
  );
  INVX1 _10205_ (
    .A( frontend_0.irq_addr_1_ ),
    .Y(_03745_)
  );
  INVX1 _10206_ (
    .A( execution_unit_0.UNUSED_inst_ad_symb ),
    .Y(_03746_)
  );
  INVX1 _10207_ (
    .A( execution_unit_0.inst_dext_15_ ),
    .Y(_03747_)
  );
  INVX1 _10208_ (
    .A( execution_unit_0.inst_dext_14_ ),
    .Y(_03748_)
  );
  INVX1 _10209_ (
    .A( execution_unit_0.inst_dext_13_ ),
    .Y(_03749_)
  );
  INVX1 _10210_ (
    .A( execution_unit_0.inst_dext_4_ ),
    .Y(_03750_)
  );
  INVX1 _10211_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .Y(_03751_)
  );
  INVX1 _10212_ (
    .A( execution_unit_0.inst_type_2_ ),
    .Y(_03752_)
  );
  INVX1 _10213_ (
    .A( execution_unit_0.inst_type_1_ ),
    .Y(_03753_)
  );
  INVX1 _10214_ (
    .A( execution_unit_0.inst_type_0_ ),
    .Y(_03754_)
  );
  INVX1 _10215_ (
    .A( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_03755_)
  );
  INVX1 _10216_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .Y(_03756_)
  );
  INVX1 _10217_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .Y(_03757_)
  );
  INVX1 _10218_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .Y(_03758_)
  );
  INVX1 _10219_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .Y(_03759_)
  );
  INVX1 _10220_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .Y(_03760_)
  );
  INVX1 _10221_ (
    .A( frontend_0.inst_dest_bin_2_ ),
    .Y(_03761_)
  );
  INVX1 _10222_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .Y(_03762_)
  );
  INVX1 _10223_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .Y(_03763_)
  );
  INVX1 _10224_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .Y(_03764_)
  );
  INVX1 _10225_ (
    .A( frontend_0.inst_src_bin_1_ ),
    .Y(_03765_)
  );
  INVX1 _10226_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .Y(_03766_)
  );
  INVX1 _10227_ (
    .A( frontend_0.inst_src_bin_0_ ),
    .Y(_03767_)
  );
  INVX1 _10228_ (
    .A( execution_unit_0.inst_as_7_ ),
    .Y(_03768_)
  );
  INVX1 _10229_ (
    .A( execution_unit_0.inst_as_4_ ),
    .Y(_03769_)
  );
  INVX1 _10230_ (
    .A( frontend_0.inst_sz_1_ ),
    .Y(_03770_)
  );
  INVX1 _10231_ (
    .A( frontend_0.exec_jmp ),
    .Y(_03771_)
  );
  INVX1 _10232_ (
    .A( frontend_0.exec_dst_wr ),
    .Y(_03772_)
  );
  INVX1 _10233_ (
    .A( frontend_0.exec_src_wr ),
    .Y(_03773_)
  );
  INVX1 _10234_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_03774_)
  );
  INVX1 _10235_ (
    .A( dbg_0.dbg_halt_cmd ),
    .Y(_03775_)
  );
  INVX1 _10236_ (
    .A( frontend_0.i_state_1_ ),
    .Y(_03776_)
  );
  INVX1 _10237_ (
    .A( frontend_0.i_state_0_ ),
    .Y(_03777_)
  );
  INVX1 _10238_ (
    .A( frontend_0.i_state_2_ ),
    .Y(_03778_)
  );
  INVX1 _10239_ (
    .A(irq_3_),
    .Y(_03779_)
  );
  INVX1 _10240_ (
    .A(irq_6_),
    .Y(_03780_)
  );
  INVX1 _10241_ (
    .A(irq_9_),
    .Y(_03781_)
  );
  INVX1 _10242_ (
    .A(irq_11_),
    .Y(_03782_)
  );
  INVX1 _10243_ (
    .A(irq_13_),
    .Y(_03783_)
  );
  INVX1 _10244_ (
    .A( execution_unit_0.gie ),
    .Y(_03784_)
  );
  INVX1 _10245_ (
    .A(1'h0),
    .Y(_03785_)
  );
  INVX1 _10246_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_03786_)
  );
  INVX1 _10247_ (
    .A( execution_unit_0.e_state_1_ ),
    .Y(_03787_)
  );
  INVX1 _10248_ (
    .A( execution_unit_0.e_state_2_ ),
    .Y(_03788_)
  );
  INVX1 _10249_ (
    .A( execution_unit_0.e_state_3_ ),
    .Y(_03789_)
  );
  INVX1 _10250_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .Y(_03790_)
  );
  INVX1 _10251_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .Y(_03791_)
  );
  INVX1 _10252_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .Y(_03792_)
  );
  INVX1 _10253_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .Y(_03793_)
  );
  INVX1 _10254_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .Y(_03794_)
  );
  INVX1 _10255_ (
    .A( execution_unit_0.pc_sw_wr ),
    .Y(_03795_)
  );
  INVX1 _10256_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_03796_)
  );
  INVX1 _10257_ (
    .A( dbg_0.UNUSED_pc_1_ ),
    .Y(_03797_)
  );
  INVX1 _10258_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .Y(_03798_)
  );
  INVX1 _10259_ (
    .A( dbg_0.UNUSED_pc_3_ ),
    .Y(_03799_)
  );
  INVX1 _10260_ (
    .A( dbg_0.UNUSED_pc_4_ ),
    .Y(_03800_)
  );
  INVX1 _10261_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .Y(_03801_)
  );
  INVX1 _10262_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .Y(_03802_)
  );
  INVX1 _10263_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .Y(_03803_)
  );
  INVX1 _10264_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .Y(_03804_)
  );
  INVX1 _10265_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .Y(_03805_)
  );
  INVX1 _10266_ (
    .A( dbg_0.UNUSED_pc_9_ ),
    .Y(_03806_)
  );
  INVX1 _10267_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .Y(_03807_)
  );
  INVX1 _10268_ (
    .A( dbg_0.UNUSED_pc_11_ ),
    .Y(_03808_)
  );
  INVX1 _10269_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .Y(_03809_)
  );
  INVX1 _10270_ (
    .A( dbg_0.UNUSED_pc_13_ ),
    .Y(_03810_)
  );
  INVX1 _10271_ (
    .A( dbg_0.UNUSED_pc_14_ ),
    .Y(_03811_)
  );
  INVX1 _10272_ (
    .A( dbg_0.UNUSED_pc_15_ ),
    .Y(_03812_)
  );
  INVX1 _10273_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .Y(_03813_)
  );
  INVX1 _10274_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .Y(_03814_)
  );
  INVX1 _10275_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03815_)
  );
  INVX1 _10276_ (
    .A( frontend_0.pmem_busy ),
    .Y(_03816_)
  );
  INVX1 _10277_ (
    .A(_06327_),
    .Y(_03254_)
  );
  NOR2X1 _10278_ (
    .A( frontend_0.i_state_1_ ),
    .B(_03777_),
    .Y(_03817_)
  );
  NAND2X1 _10279_ (
    .A(_03776_),
    .B( frontend_0.i_state_0_ ),
    .Y(_03818_)
  );
  NOR2X1 _10280_ (
    .A(_03778_),
    .B(_03818_),
    .Y(_03819_)
  );
  NAND2X1 _10281_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03817_),
    .Y(_03820_)
  );
  OR2X1 _10282_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03821_)
  );
  NAND2X1 _10283_ (
    .A( execution_unit_0.e_state_2_ ),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_03822_)
  );
  OAI21X1 _10284_ (
    .A(_03821_),
    .B(_03822_),
    .C( frontend_0.exec_jmp ),
    .Y(_03823_)
  );
  INVX1 _10285_ (
    .A(_03823_),
    .Y(_03824_)
  );
  NAND2X1 _10286_ (
    .A(_03788_),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_03825_)
  );
  OR2X1 _10287_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03787_),
    .Y(_03826_)
  );
  NOR2X1 _10288_ (
    .A(_03825_),
    .B(_03826_),
    .Y(_03827_)
  );
  OR2X1 _10289_ (
    .A(_03825_),
    .B(_03826_),
    .Y(_03828_)
  );
  AND2X1 _10290_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03829_)
  );
  NAND2X1 _10291_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03830_)
  );
  NAND2X1 _10292_ (
    .A( execution_unit_0.e_state_2_ ),
    .B(_03789_),
    .Y(_03831_)
  );
  NOR3X1 _10293_ (
    .A(_03788_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_03830_),
    .Y(_03832_)
  );
  NAND3X1 _10294_ (
    .A( execution_unit_0.e_state_2_ ),
    .B(_03789_),
    .C(_03829_),
    .Y(_03833_)
  );
  NOR3X1 _10295_ (
    .A( execution_unit_0.e_state_2_ ),
    .B(_03789_),
    .C(_03830_),
    .Y(_03834_)
  );
  NAND3X1 _10296_ (
    .A(_03788_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_03829_),
    .Y(_03835_)
  );
  MUX2X1 _10297_ (
    .A(_03832_),
    .B(_03834_),
    .S( frontend_0.exec_src_wr ),
    .Y(_03836_)
  );
  MUX2X1 _10298_ (
    .A(_03828_),
    .B(_03836_),
    .S( frontend_0.exec_dst_wr ),
    .Y(_03837_)
  );
  OAI21X1 _10299_ (
    .A( frontend_0.exec_jmp ),
    .B(_03837_),
    .C(_03823_),
    .Y(_03838_)
  );
  INVX1 _10300_ (
    .A(_03838_),
    .Y( execution_unit_0.exec_done )
  );
  NOR2X1 _10301_ (
    .A(irq_3_),
    .B(irq_2_),
    .Y(_03839_)
  );
  NOR2X1 _10302_ (
    .A(irq_9_),
    .B(irq_8_),
    .Y(_03840_)
  );
  INVX1 _10303_ (
    .A(_03840_),
    .Y(_03841_)
  );
  NOR2X1 _10304_ (
    .A(irq_13_),
    .B(irq_12_),
    .Y(_03842_)
  );
  NOR2X1 _10305_ (
    .A(irq_7_),
    .B(irq_6_),
    .Y(_03843_)
  );
  OR2X1 _10306_ (
    .A(irq_7_),
    .B(irq_6_),
    .Y(_03844_)
  );
  NAND2X1 _10307_ (
    .A(_03840_),
    .B(_03842_),
    .Y(_03845_)
  );
  NAND2X1 _10308_ (
    .A(_03839_),
    .B(_03843_),
    .Y(_03846_)
  );
  OR2X1 _10309_ (
    .A(irq_10_),
    .B( frontend_0.wdt_irq ),
    .Y(_03847_)
  );
  NOR3X1 _10310_ (
    .A(irq_11_),
    .B(irq_10_),
    .C( frontend_0.wdt_irq ),
    .Y(_03848_)
  );
  NOR2X1 _10311_ (
    .A(irq_0_),
    .B(irq_5_),
    .Y(_03849_)
  );
  NOR2X1 _10312_ (
    .A(irq_1_),
    .B(irq_4_),
    .Y(_03850_)
  );
  NAND3X1 _10313_ (
    .A(_03848_),
    .B(_03849_),
    .C(_03850_),
    .Y(_03851_)
  );
  NOR3X1 _10314_ (
    .A(_03845_),
    .B(_03846_),
    .C(_03851_),
    .Y(_03852_)
  );
  OAI21X1 _10315_ (
    .A(_03784_),
    .B(_03852_),
    .C(_03785_),
    .Y(_03853_)
  );
  AND2X1 _10316_ (
    .A(_03775_),
    .B(cpu_en),
    .Y(_03854_)
  );
  NAND2X1 _10317_ (
    .A(_03775_),
    .B(cpu_en),
    .Y(_03855_)
  );
  NOR2X1 _10318_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_03855_),
    .Y(_03856_)
  );
  AND2X1 _10319_ (
    .A(_03853_),
    .B(_03856_),
    .Y(_03857_)
  );
  NAND2X1 _10320_ (
    .A(_03853_),
    .B(_03856_),
    .Y(_03858_)
  );
  AOI21X1 _10321_ (
    .A(_03820_),
    .B(_03838_),
    .C(_03858_),
    .Y(_03859_)
  );
  OAI21X1 _10322_ (
    .A(_03819_),
    .B( execution_unit_0.exec_done ),
    .C(_03857_),
    .Y(_03860_)
  );
  NAND2X1 _10323_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03860_),
    .Y(_03861_)
  );
  NOR2X1 _10324_ (
    .A(irq_7_),
    .B(_03780_),
    .Y(_03862_)
  );
  AOI21X1 _10325_ (
    .A(_03783_),
    .B(irq_12_),
    .C(1'h0),
    .Y(_03863_)
  );
  NAND3X1 _10326_ (
    .A(_03841_),
    .B(_03848_),
    .C(_03863_),
    .Y(_03864_)
  );
  OAI21X1 _10327_ (
    .A(1'h0),
    .B(_03842_),
    .C(_03864_),
    .Y(_03865_)
  );
  INVX1 _10328_ (
    .A(_03865_),
    .Y(_03866_)
  );
  AND2X1 _10329_ (
    .A(_03785_),
    .B(_03842_),
    .Y(_03867_)
  );
  NAND2X1 _10330_ (
    .A(_03840_),
    .B(_03848_),
    .Y(_03868_)
  );
  NAND2X1 _10331_ (
    .A(_03867_),
    .B(_03868_),
    .Y(_03869_)
  );
  AND2X1 _10332_ (
    .A(_03866_),
    .B(_03869_),
    .Y(_03870_)
  );
  AOI21X1 _10333_ (
    .A(_03781_),
    .B(irq_8_),
    .C(_03847_),
    .Y(_03871_)
  );
  NAND2X1 _10334_ (
    .A(_03782_),
    .B(_03867_),
    .Y(_03872_)
  );
  OAI21X1 _10335_ (
    .A(_03871_),
    .B(_03872_),
    .C(_03863_),
    .Y(_03873_)
  );
  INVX1 _10336_ (
    .A(_03873_),
    .Y(_03874_)
  );
  NAND2X1 _10337_ (
    .A(_03870_),
    .B(_03874_),
    .Y(_03875_)
  );
  OAI21X1 _10338_ (
    .A(irq_7_),
    .B(_03780_),
    .C(irq_4_),
    .Y(_03876_)
  );
  AOI21X1 _10339_ (
    .A(_03862_),
    .B(_03870_),
    .C(_03873_),
    .Y(_03877_)
  );
  NOR2X1 _10340_ (
    .A(_03875_),
    .B(_03876_),
    .Y(_03878_)
  );
  NOR2X1 _10341_ (
    .A(irq_5_),
    .B(_03844_),
    .Y(_03879_)
  );
  NOR2X1 _10342_ (
    .A(_03875_),
    .B(_03879_),
    .Y(_03880_)
  );
  NOR2X1 _10343_ (
    .A(_03878_),
    .B(_03880_),
    .Y(_03881_)
  );
  NAND2X1 _10344_ (
    .A(_03878_),
    .B(_03879_),
    .Y(_03882_)
  );
  NAND2X1 _10345_ (
    .A(_03866_),
    .B(_03882_),
    .Y(_03883_)
  );
  NOR2X1 _10346_ (
    .A(_03844_),
    .B(_03875_),
    .Y(_03884_)
  );
  AOI21X1 _10347_ (
    .A(irq_5_),
    .B(_03884_),
    .C(_03883_),
    .Y(_03885_)
  );
  INVX1 _10348_ (
    .A(_03885_),
    .Y(_03886_)
  );
  AND2X1 _10349_ (
    .A(_03869_),
    .B(_03881_),
    .Y(_03887_)
  );
  NAND3X1 _10350_ (
    .A(_03877_),
    .B(_03885_),
    .C(_03887_),
    .Y(_03888_)
  );
  OAI21X1 _10351_ (
    .A(_03839_),
    .B(_03888_),
    .C(_03881_),
    .Y(_03889_)
  );
  NAND2X1 _10352_ (
    .A(_03779_),
    .B(irq_2_),
    .Y(_03890_)
  );
  AND2X1 _10353_ (
    .A(_03877_),
    .B(_03882_),
    .Y(_03891_)
  );
  OAI21X1 _10354_ (
    .A(_03888_),
    .B(_03890_),
    .C(_03891_),
    .Y(_03892_)
  );
  OAI21X1 _10355_ (
    .A(_03839_),
    .B(_03888_),
    .C(_03869_),
    .Y(_03893_)
  );
  NOR2X1 _10356_ (
    .A(_03892_),
    .B(_03893_),
    .Y(_03894_)
  );
  NAND2X1 _10357_ (
    .A(irq_1_),
    .B(_03885_),
    .Y(_03895_)
  );
  NOR2X1 _10358_ (
    .A(_03889_),
    .B(_03895_),
    .Y(_03896_)
  );
  AND2X1 _10359_ (
    .A(_03894_),
    .B(_03896_),
    .Y(_03897_)
  );
  NAND2X1 _10360_ (
    .A(irq_0_),
    .B(_03885_),
    .Y(_03898_)
  );
  NOR2X1 _10361_ (
    .A(_03889_),
    .B(_03898_),
    .Y(_03899_)
  );
  NAND2X1 _10362_ (
    .A(_03894_),
    .B(_03899_),
    .Y(_03900_)
  );
  OAI21X1 _10363_ (
    .A(_03896_),
    .B(_03900_),
    .C(_03859_),
    .Y(_03901_)
  );
  OR2X1 _10364_ (
    .A(_03897_),
    .B(_03901_),
    .Y(_03902_)
  );
  OAI21X1 _10365_ (
    .A(_03889_),
    .B(_03902_),
    .C(_03861_),
    .Y(_03454_)
  );
  OAI22X1 _10366_ (
    .A(_03743_),
    .B(_03859_),
    .C(_03893_),
    .D(_03902_),
    .Y(_03453_)
  );
  OAI22X1 _10367_ (
    .A(_03744_),
    .B(_03859_),
    .C(_03886_),
    .D(_03902_),
    .Y(_03452_)
  );
  OAI22X1 _10368_ (
    .A(_03745_),
    .B(_03859_),
    .C(_03892_),
    .D(_03901_),
    .Y(_03451_)
  );
  AND2X1 _10369_ (
    .A( execution_unit_0.inst_irq_rst ),
    .B(_03838_),
    .Y(_03450_)
  );
  NAND2X1 _10370_ (
    .A( frontend_0.i_state_1_ ),
    .B(_03778_),
    .Y(_03903_)
  );
  NOR2X1 _10371_ (
    .A( frontend_0.i_state_0_ ),
    .B(_03903_),
    .Y(_03904_)
  );
  INVX1 _10372_ (
    .A(_03904_),
    .Y(_03905_)
  );
  NAND2X1 _10373_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03787_),
    .Y(_03906_)
  );
  OR2X1 _10374_ (
    .A(_03822_),
    .B(_03906_),
    .Y(_03907_)
  );
  OAI21X1 _10375_ (
    .A(_03822_),
    .B(_03906_),
    .C(_03838_),
    .Y(_03908_)
  );
  NAND2X1 _10376_ (
    .A(_03904_),
    .B(_03908_),
    .Y(_03909_)
  );
  INVX1 _10377_ (
    .A(_03909_),
    .Y( dbg_0.decode_noirq )
  );
  NOR2X1 _10378_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .Y(_03910_)
  );
  NAND2X1 _10379_ (
    .A(_03860_),
    .B(_03909_),
    .Y(_03911_)
  );
  NAND2X1 _10380_ (
    .A( execution_unit_0.inst_ad_6_ ),
    .B(_03910_),
    .Y(_03912_)
  );
  NOR2X1 _10381_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .Y(_03913_)
  );
  OR2X1 _10382_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .Y(_03914_)
  );
  NAND2X1 _10383_ (
    .A(_03860_),
    .B( dbg_0.decode_noirq ),
    .Y(_03915_)
  );
  INVX1 _10384_ (
    .A(_03915_),
    .Y(_03916_)
  );
  NOR2X1 _10385_ (
    .A(_03859_),
    .B(_03913_),
    .Y(_03917_)
  );
  OAI21X1 _10386_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .C(_03916_),
    .Y(_03918_)
  );
  NOR2X1 _10387_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B( dbg_0.fe_mdb_in_2_ ),
    .Y(_03919_)
  );
  OR2X1 _10388_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B( dbg_0.fe_mdb_in_2_ ),
    .Y(_03920_)
  );
  NOR2X1 _10389_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03920_),
    .Y(_03921_)
  );
  NAND3X1 _10390_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B( dbg_0.fe_mdb_in_7_ ),
    .C(_03921_),
    .Y(_03922_)
  );
  OAI21X1 _10391_ (
    .A(_03918_),
    .B(_03922_),
    .C(_03912_),
    .Y(_03449_)
  );
  AND2X1 _10392_ (
    .A(_03762_),
    .B(_03921_),
    .Y(_03923_)
  );
  AND2X1 _10393_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03917_),
    .Y(_03924_)
  );
  NAND2X1 _10394_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03917_),
    .Y(_03925_)
  );
  OAI21X1 _10395_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03924_),
    .Y(_03926_)
  );
  NAND3X1 _10396_ (
    .A(_03911_),
    .B(_03923_),
    .C(_03924_),
    .Y(_03927_)
  );
  OAI21X1 _10397_ (
    .A(_03746_),
    .B(_03911_),
    .C(_03927_),
    .Y(_03448_)
  );
  NAND2X1 _10398_ (
    .A( execution_unit_0.UNUSED_inst_ad_idx ),
    .B(_03910_),
    .Y(_03928_)
  );
  OAI21X1 _10399_ (
    .A(_03921_),
    .B(_03926_),
    .C(_03928_),
    .Y(_03447_)
  );
  NAND2X1 _10400_ (
    .A( execution_unit_0.inst_ad_0_ ),
    .B(_03910_),
    .Y(_03929_)
  );
  NOR2X1 _10401_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03918_),
    .Y(_03930_)
  );
  OAI21X1 _10402_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03918_),
    .C(_03929_),
    .Y(_03446_)
  );
  NOR3X1 _10403_ (
    .A(_03791_),
    .B(_03859_),
    .C(_03914_),
    .Y(_03931_)
  );
  NAND3X1 _10404_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03860_),
    .C(_03913_),
    .Y(_03932_)
  );
  NOR2X1 _10405_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03914_),
    .Y(_03933_)
  );
  NAND2X1 _10406_ (
    .A(_03791_),
    .B(_03913_),
    .Y(_03934_)
  );
  NAND2X1 _10407_ (
    .A(_03860_),
    .B(_03933_),
    .Y(_03935_)
  );
  NOR2X1 _10408_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( dbg_0.fe_mdb_in_10_ ),
    .Y(_03936_)
  );
  OR2X1 _10409_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( dbg_0.fe_mdb_in_10_ ),
    .Y(_03937_)
  );
  AOI21X1 _10410_ (
    .A(_03860_),
    .B(_03933_),
    .C(_03937_),
    .Y(_03938_)
  );
  OAI21X1 _10411_ (
    .A(_03859_),
    .B(_03934_),
    .C(_03936_),
    .Y(_03939_)
  );
  NOR3X1 _10412_ (
    .A(_03859_),
    .B(_03920_),
    .C(_03934_),
    .Y(_03940_)
  );
  NAND3X1 _10413_ (
    .A(_03860_),
    .B(_03919_),
    .C(_03933_),
    .Y(_03941_)
  );
  NOR3X1 _10414_ (
    .A(_03762_),
    .B(_03859_),
    .C(_03934_),
    .Y(_03942_)
  );
  NAND3X1 _10415_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B(_03860_),
    .C(_03933_),
    .Y(_03943_)
  );
  AOI21X1 _10416_ (
    .A(_03860_),
    .B(_03933_),
    .C(_03764_),
    .Y(_03944_)
  );
  OAI21X1 _10417_ (
    .A(_03859_),
    .B(_03934_),
    .C( dbg_0.fe_mdb_in_9_ ),
    .Y(_03945_)
  );
  NOR2X1 _10418_ (
    .A(_03942_),
    .B(_03944_),
    .Y(_03946_)
  );
  OAI21X1 _10419_ (
    .A(_03762_),
    .B(_03935_),
    .C(_03945_),
    .Y(_03947_)
  );
  AOI22X1 _10420_ (
    .A(_03939_),
    .B(_03941_),
    .C(_03943_),
    .D(_03945_),
    .Y(_03948_)
  );
  OAI22X1 _10421_ (
    .A(_03938_),
    .B(_03940_),
    .C(_03942_),
    .D(_03944_),
    .Y(_03949_)
  );
  AOI21X1 _10422_ (
    .A(_03860_),
    .B(_03933_),
    .C( dbg_0.fe_mdb_in_8_ ),
    .Y(_03950_)
  );
  OAI21X1 _10423_ (
    .A(_03859_),
    .B(_03934_),
    .C(_03766_),
    .Y(_03951_)
  );
  NOR3X1 _10424_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03859_),
    .C(_03934_),
    .Y(_03952_)
  );
  NAND3X1 _10425_ (
    .A(_03751_),
    .B(_03860_),
    .C(_03933_),
    .Y(_03953_)
  );
  NOR2X1 _10426_ (
    .A(_03950_),
    .B(_03952_),
    .Y(_03954_)
  );
  AND2X1 _10427_ (
    .A(_03948_),
    .B(_03954_),
    .Y(_03955_)
  );
  NAND2X1 _10428_ (
    .A(_03932_),
    .B(_03955_),
    .Y(_03956_)
  );
  AOI22X1 _10429_ (
    .A(_03939_),
    .B(_03941_),
    .C(_03951_),
    .D(_03953_),
    .Y(_03957_)
  );
  OAI22X1 _10430_ (
    .A(_03938_),
    .B(_03940_),
    .C(_03950_),
    .D(_03952_),
    .Y(_03958_)
  );
  OAI21X1 _10431_ (
    .A(_03950_),
    .B(_03952_),
    .C(_03948_),
    .Y(_03959_)
  );
  NAND2X1 _10432_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03932_),
    .Y(_03960_)
  );
  OAI21X1 _10433_ (
    .A(_03959_),
    .B(_03960_),
    .C(_03956_),
    .Y(_03961_)
  );
  AND2X1 _10434_ (
    .A(_03911_),
    .B(_03961_),
    .Y(_03962_)
  );
  OAI21X1 _10435_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03961_),
    .Y(_03963_)
  );
  NOR2X1 _10436_ (
    .A(_03909_),
    .B(_03932_),
    .Y(_03964_)
  );
  NAND2X1 _10437_ (
    .A( dbg_0.decode_noirq ),
    .B(_03931_),
    .Y(_03965_)
  );
  NOR2X1 _10438_ (
    .A(_03764_),
    .B(_03965_),
    .Y(_03966_)
  );
  NAND2X1 _10439_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03964_),
    .Y(_03967_)
  );
  NOR2X1 _10440_ (
    .A(_03777_),
    .B(_03903_),
    .Y(_03968_)
  );
  OR2X1 _10441_ (
    .A(_03777_),
    .B(_03903_),
    .Y(_03969_)
  );
  NOR2X1 _10442_ (
    .A( frontend_0.i_state_1_ ),
    .B( frontend_0.i_state_0_ ),
    .Y(_03970_)
  );
  NAND2X1 _10443_ (
    .A(_03776_),
    .B(_03777_),
    .Y(_03971_)
  );
  NAND2X1 _10444_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03970_),
    .Y(_03972_)
  );
  AOI21X1 _10445_ (
    .A(_03770_),
    .B( frontend_0.inst_sz_0_ ),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03973_)
  );
  INVX1 _10446_ (
    .A(_03973_),
    .Y(_03974_)
  );
  NAND2X1 _10447_ (
    .A(_03968_),
    .B(_03974_),
    .Y(_03975_)
  );
  OAI21X1 _10448_ (
    .A( execution_unit_0.inst_as_4_ ),
    .B(_03975_),
    .C(_03972_),
    .Y(_03976_)
  );
  NAND2X1 _10449_ (
    .A( execution_unit_0.UNUSED_inst_ad_symb ),
    .B(_03976_),
    .Y(_03977_)
  );
  AOI22X1 _10450_ (
    .A( execution_unit_0.inst_as_4_ ),
    .B(_03968_),
    .C(_03976_),
    .D( execution_unit_0.UNUSED_inst_ad_symb ),
    .Y(_03978_)
  );
  OAI21X1 _10451_ (
    .A(_03769_),
    .B(_03969_),
    .C(_03977_),
    .Y(_03979_)
  );
  XNOR2X1 _10452_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03978_),
    .Y(_03980_)
  );
  XNOR2X1 _10453_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B(_03978_),
    .Y(_03981_)
  );
  AND2X1 _10454_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B(_03979_),
    .Y(_03982_)
  );
  NAND2X1 _10455_ (
    .A(_03793_),
    .B(_03919_),
    .Y(_03983_)
  );
  NOR2X1 _10456_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B( dbg_0.fe_mdb_in_8_ ),
    .Y(_03984_)
  );
  NOR2X1 _10457_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_03985_)
  );
  NAND3X1 _10458_ (
    .A(_03803_),
    .B(_03984_),
    .C(_03985_),
    .Y(_03986_)
  );
  OR2X1 _10459_ (
    .A(_03983_),
    .B(_03986_),
    .Y(_03987_)
  );
  NOR2X1 _10460_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03987_),
    .Y(_03988_)
  );
  NAND3X1 _10461_ (
    .A(_03762_),
    .B(_03793_),
    .C(_03919_),
    .Y(_03989_)
  );
  OR2X1 _10462_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03989_),
    .Y(_03990_)
  );
  NOR2X1 _10463_ (
    .A(_03978_),
    .B(_03988_),
    .Y(_03991_)
  );
  NOR2X1 _10464_ (
    .A(_03982_),
    .B(_03991_),
    .Y(_03992_)
  );
  OAI21X1 _10465_ (
    .A(_03982_),
    .B(_03991_),
    .C(_03981_),
    .Y(_03993_)
  );
  INVX1 _10466_ (
    .A(_03993_),
    .Y(_03994_)
  );
  AOI21X1 _10467_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B(_03979_),
    .C(_03994_),
    .Y(_03995_)
  );
  XNOR2X1 _10468_ (
    .A(_03756_),
    .B(_03978_),
    .Y(_03996_)
  );
  OAI21X1 _10469_ (
    .A(_03756_),
    .B(_03978_),
    .C(_03995_),
    .Y(_03997_)
  );
  NAND2X1 _10470_ (
    .A(_03980_),
    .B(_03997_),
    .Y(_03998_)
  );
  OAI21X1 _10471_ (
    .A(_03791_),
    .B(_03978_),
    .C(_03998_),
    .Y(_03999_)
  );
  INVX1 _10472_ (
    .A(_03999_),
    .Y(_04000_)
  );
  OAI21X1 _10473_ (
    .A(_03790_),
    .B(_03978_),
    .C(_04000_),
    .Y(_04001_)
  );
  XNOR2X1 _10474_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03978_),
    .Y(_04002_)
  );
  XOR2X1 _10475_ (
    .A(_04001_),
    .B(_04002_),
    .Y(_04003_)
  );
  OAI21X1 _10476_ (
    .A(_03966_),
    .B(_04003_),
    .C(_03963_),
    .Y(_04004_)
  );
  NOR2X1 _10477_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B( execution_unit_0.inst_as_5_ ),
    .Y(_04005_)
  );
  NOR2X1 _10478_ (
    .A( execution_unit_0.inst_as_4_ ),
    .B( execution_unit_0.inst_as_1_ ),
    .Y(_04006_)
  );
  NAND2X1 _10479_ (
    .A(_04005_),
    .B(_04006_),
    .Y(_04007_)
  );
  NAND2X1 _10480_ (
    .A(_03968_),
    .B(_04007_),
    .Y(_04008_)
  );
  INVX1 _10481_ (
    .A(_04008_),
    .Y(_04009_)
  );
  OAI21X1 _10482_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04008_),
    .Y(_04010_)
  );
  NOR2X1 _10483_ (
    .A(_03962_),
    .B(_04010_),
    .Y(_04011_)
  );
  OR2X1 _10484_ (
    .A(_03962_),
    .B(_04010_),
    .Y(_04012_)
  );
  NAND2X1 _10485_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03932_),
    .Y(_04013_)
  );
  NOR3X1 _10486_ (
    .A(_03792_),
    .B(_03793_),
    .C(_03931_),
    .Y(_04014_)
  );
  NAND3X1 _10487_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B( dbg_0.fe_mdb_in_4_ ),
    .C(_03932_),
    .Y(_04015_)
  );
  NAND2X1 _10488_ (
    .A(_03948_),
    .B(_04014_),
    .Y(_04016_)
  );
  NOR2X1 _10489_ (
    .A(_03963_),
    .B(_04016_),
    .Y(_04017_)
  );
  AOI21X1 _10490_ (
    .A(_03954_),
    .B(_04017_),
    .C(_04011_),
    .Y(_04018_)
  );
  NOR2X1 _10491_ (
    .A( execution_unit_0.inst_sext_15_ ),
    .B(_04012_),
    .Y(_04019_)
  );
  AOI21X1 _10492_ (
    .A(_04004_),
    .B(_04018_),
    .C(_04019_),
    .Y(_03445_)
  );
  XNOR2X1 _10493_ (
    .A(_03790_),
    .B(_03978_),
    .Y(_04020_)
  );
  XNOR2X1 _10494_ (
    .A(_03999_),
    .B(_04020_),
    .Y(_04021_)
  );
  OAI21X1 _10495_ (
    .A(_03966_),
    .B(_04021_),
    .C(_03963_),
    .Y(_04022_)
  );
  NOR2X1 _10496_ (
    .A( execution_unit_0.inst_sext_14_ ),
    .B(_04012_),
    .Y(_04023_)
  );
  AOI21X1 _10497_ (
    .A(_04018_),
    .B(_04022_),
    .C(_04023_),
    .Y(_03444_)
  );
  XOR2X1 _10498_ (
    .A(_03980_),
    .B(_03997_),
    .Y(_04024_)
  );
  AOI21X1 _10499_ (
    .A(_03965_),
    .B(_04024_),
    .C(_03966_),
    .Y(_04025_)
  );
  OAI21X1 _10500_ (
    .A(_03962_),
    .B(_04025_),
    .C(_04018_),
    .Y(_04026_)
  );
  OAI21X1 _10501_ (
    .A( execution_unit_0.inst_sext_13_ ),
    .B(_04012_),
    .C(_04026_),
    .Y(_04027_)
  );
  INVX1 _10502_ (
    .A(_04027_),
    .Y(_03443_)
  );
  XNOR2X1 _10503_ (
    .A(_03995_),
    .B(_03996_),
    .Y(_04028_)
  );
  OAI21X1 _10504_ (
    .A(_03964_),
    .B(_04028_),
    .C(_03967_),
    .Y(_04029_)
  );
  NAND2X1 _10505_ (
    .A(_03963_),
    .B(_04029_),
    .Y(_04030_)
  );
  NOR2X1 _10506_ (
    .A( execution_unit_0.inst_sext_12_ ),
    .B(_04012_),
    .Y(_04031_)
  );
  AOI21X1 _10507_ (
    .A(_04018_),
    .B(_04030_),
    .C(_04031_),
    .Y(_03442_)
  );
  XOR2X1 _10508_ (
    .A(_03981_),
    .B(_03992_),
    .Y(_04032_)
  );
  OAI21X1 _10509_ (
    .A(_03964_),
    .B(_04032_),
    .C(_03967_),
    .Y(_04033_)
  );
  NAND2X1 _10510_ (
    .A(_03963_),
    .B(_04033_),
    .Y(_04034_)
  );
  NOR2X1 _10511_ (
    .A( execution_unit_0.inst_sext_11_ ),
    .B(_04012_),
    .Y(_04035_)
  );
  AOI21X1 _10512_ (
    .A(_04018_),
    .B(_04034_),
    .C(_04035_),
    .Y(_03441_)
  );
  NOR2X1 _10513_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B(_03979_),
    .Y(_04036_)
  );
  NOR2X1 _10514_ (
    .A(_03982_),
    .B(_04036_),
    .Y(_04037_)
  );
  XNOR2X1 _10515_ (
    .A(_03991_),
    .B(_04037_),
    .Y(_04038_)
  );
  OAI21X1 _10516_ (
    .A(_03964_),
    .B(_04038_),
    .C(_03967_),
    .Y(_04039_)
  );
  NAND2X1 _10517_ (
    .A(_03963_),
    .B(_04039_),
    .Y(_04040_)
  );
  NOR2X1 _10518_ (
    .A( execution_unit_0.inst_sext_10_ ),
    .B(_04012_),
    .Y(_04041_)
  );
  AOI21X1 _10519_ (
    .A(_04018_),
    .B(_04040_),
    .C(_04041_),
    .Y(_03440_)
  );
  NAND2X1 _10520_ (
    .A(_03762_),
    .B(_03979_),
    .Y(_04042_)
  );
  NOR2X1 _10521_ (
    .A(_03978_),
    .B(_03989_),
    .Y(_04043_)
  );
  NOR2X1 _10522_ (
    .A(_03978_),
    .B(_03990_),
    .Y(_04044_)
  );
  NAND2X1 _10523_ (
    .A(_03803_),
    .B(_04044_),
    .Y(_04045_)
  );
  OR2X1 _10524_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_04045_),
    .Y(_04046_)
  );
  NOR2X1 _10525_ (
    .A(_03978_),
    .B(_03987_),
    .Y(_04047_)
  );
  XNOR2X1 _10526_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_04047_),
    .Y(_04048_)
  );
  OAI21X1 _10527_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04048_),
    .Y(_04049_)
  );
  OAI21X1 _10528_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03965_),
    .C(_04049_),
    .Y(_04050_)
  );
  OAI21X1 _10529_ (
    .A(_03962_),
    .B(_04050_),
    .C(_04018_),
    .Y(_04051_)
  );
  OAI21X1 _10530_ (
    .A( execution_unit_0.inst_sext_9_ ),
    .B(_04012_),
    .C(_04051_),
    .Y(_04052_)
  );
  INVX1 _10531_ (
    .A(_04052_),
    .Y(_03439_)
  );
  XNOR2X1 _10532_ (
    .A(_03766_),
    .B(_04046_),
    .Y(_04053_)
  );
  OAI21X1 _10533_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04053_),
    .Y(_04054_)
  );
  OAI21X1 _10534_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03965_),
    .C(_04054_),
    .Y(_04055_)
  );
  OAI21X1 _10535_ (
    .A(_03962_),
    .B(_04055_),
    .C(_04018_),
    .Y(_04056_)
  );
  OAI21X1 _10536_ (
    .A( execution_unit_0.inst_sext_8_ ),
    .B(_04012_),
    .C(_04056_),
    .Y(_04057_)
  );
  INVX1 _10537_ (
    .A(_04057_),
    .Y(_03438_)
  );
  XNOR2X1 _10538_ (
    .A(_03794_),
    .B(_04045_),
    .Y(_04058_)
  );
  OAI21X1 _10539_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04058_),
    .Y(_04059_)
  );
  OAI21X1 _10540_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03965_),
    .C(_04059_),
    .Y(_04060_)
  );
  OAI21X1 _10541_ (
    .A(_03962_),
    .B(_04060_),
    .C(_04018_),
    .Y(_04061_)
  );
  OAI21X1 _10542_ (
    .A( execution_unit_0.inst_sext_7_ ),
    .B(_04012_),
    .C(_04061_),
    .Y(_04062_)
  );
  INVX1 _10543_ (
    .A(_04062_),
    .Y(_03437_)
  );
  OAI21X1 _10544_ (
    .A(_03978_),
    .B(_03990_),
    .C( dbg_0.fe_mdb_in_6_ ),
    .Y(_04063_)
  );
  AND2X1 _10545_ (
    .A(_04045_),
    .B(_04063_),
    .Y(_04064_)
  );
  OAI21X1 _10546_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04064_),
    .Y(_04065_)
  );
  OAI21X1 _10547_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03965_),
    .C(_04065_),
    .Y(_04066_)
  );
  OAI21X1 _10548_ (
    .A(_03962_),
    .B(_04066_),
    .C(_04018_),
    .Y(_04067_)
  );
  OAI21X1 _10549_ (
    .A( execution_unit_0.inst_sext_6_ ),
    .B(_04012_),
    .C(_04067_),
    .Y(_04068_)
  );
  INVX1 _10550_ (
    .A(_04068_),
    .Y(_03436_)
  );
  NOR2X1 _10551_ (
    .A(_03792_),
    .B(_04043_),
    .Y(_04069_)
  );
  NOR2X1 _10552_ (
    .A(_04044_),
    .B(_04069_),
    .Y(_04070_)
  );
  OAI21X1 _10553_ (
    .A(_03909_),
    .B(_03932_),
    .C(_04070_),
    .Y(_04071_)
  );
  OAI21X1 _10554_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03965_),
    .C(_04071_),
    .Y(_04072_)
  );
  OAI21X1 _10555_ (
    .A(_03962_),
    .B(_04072_),
    .C(_04018_),
    .Y(_04073_)
  );
  OAI21X1 _10556_ (
    .A( execution_unit_0.inst_sext_5_ ),
    .B(_04012_),
    .C(_04073_),
    .Y(_04074_)
  );
  INVX1 _10557_ (
    .A(_04074_),
    .Y(_03435_)
  );
  NAND2X1 _10558_ (
    .A(_03759_),
    .B(_03964_),
    .Y(_04075_)
  );
  NOR2X1 _10559_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_04042_),
    .Y(_04076_)
  );
  OAI21X1 _10560_ (
    .A(_03920_),
    .B(_04042_),
    .C( dbg_0.fe_mdb_in_4_ ),
    .Y(_04077_)
  );
  OAI21X1 _10561_ (
    .A(_03978_),
    .B(_03989_),
    .C(_04077_),
    .Y(_04078_)
  );
  OAI21X1 _10562_ (
    .A(_03964_),
    .B(_04078_),
    .C(_04075_),
    .Y(_04079_)
  );
  OAI21X1 _10563_ (
    .A(_03962_),
    .B(_04079_),
    .C(_04018_),
    .Y(_04080_)
  );
  OAI21X1 _10564_ (
    .A( execution_unit_0.inst_sext_4_ ),
    .B(_04012_),
    .C(_04080_),
    .Y(_04081_)
  );
  INVX1 _10565_ (
    .A(_04081_),
    .Y(_03434_)
  );
  XNOR2X1 _10566_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B(_04076_),
    .Y(_04082_)
  );
  NOR2X1 _10567_ (
    .A(_03964_),
    .B(_04082_),
    .Y(_04083_)
  );
  AOI21X1 _10568_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_03964_),
    .C(_04083_),
    .Y(_04084_)
  );
  OAI21X1 _10569_ (
    .A(_03962_),
    .B(_04084_),
    .C(_04012_),
    .Y(_04085_)
  );
  OAI22X1 _10570_ (
    .A( execution_unit_0.inst_sext_3_ ),
    .B(_04012_),
    .C(_04017_),
    .D(_04085_),
    .Y(_04086_)
  );
  INVX1 _10571_ (
    .A(_04086_),
    .Y(_03433_)
  );
  NOR2X1 _10572_ (
    .A( execution_unit_0.inst_sext_2_ ),
    .B(_04012_),
    .Y(_04087_)
  );
  XOR2X1 _10573_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_04042_),
    .Y(_04088_)
  );
  MUX2X1 _10574_ (
    .A(_03762_),
    .B(_04088_),
    .S(_03964_),
    .Y(_04089_)
  );
  NOR3X1 _10575_ (
    .A(_03792_),
    .B( dbg_0.fe_mdb_in_4_ ),
    .C(_03931_),
    .Y(_04090_)
  );
  NAND3X1 _10576_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03793_),
    .C(_03932_),
    .Y(_04091_)
  );
  OAI21X1 _10577_ (
    .A(_03959_),
    .B(_04091_),
    .C(_03962_),
    .Y(_04092_)
  );
  OAI21X1 _10578_ (
    .A(_03962_),
    .B(_04089_),
    .C(_04092_),
    .Y(_04093_)
  );
  AOI21X1 _10579_ (
    .A(_04018_),
    .B(_04093_),
    .C(_04087_),
    .Y(_03432_)
  );
  NAND2X1 _10580_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03964_),
    .Y(_04094_)
  );
  XNOR2X1 _10581_ (
    .A(_03762_),
    .B(_03978_),
    .Y(_04095_)
  );
  OAI21X1 _10582_ (
    .A(_03964_),
    .B(_04095_),
    .C(_04094_),
    .Y(_04096_)
  );
  NOR2X1 _10583_ (
    .A(_03910_),
    .B(_03960_),
    .Y(_04097_)
  );
  AOI22X1 _10584_ (
    .A(_03963_),
    .B(_04096_),
    .C(_04097_),
    .D(_03955_),
    .Y(_04098_)
  );
  NAND2X1 _10585_ (
    .A( execution_unit_0.inst_sext_1_ ),
    .B(_04011_),
    .Y(_04099_)
  );
  OAI21X1 _10586_ (
    .A(_04011_),
    .B(_04098_),
    .C(_04099_),
    .Y(_03431_)
  );
  NOR2X1 _10587_ (
    .A(_03751_),
    .B(_03964_),
    .Y(_04100_)
  );
  NOR2X1 _10588_ (
    .A(_03793_),
    .B(_03956_),
    .Y(_04101_)
  );
  AOI22X1 _10589_ (
    .A(_03963_),
    .B(_04100_),
    .C(_04101_),
    .D(_03911_),
    .Y(_04102_)
  );
  NAND2X1 _10590_ (
    .A( execution_unit_0.inst_sext_0_ ),
    .B(_04011_),
    .Y(_04103_)
  );
  OAI21X1 _10591_ (
    .A(_04011_),
    .B(_04102_),
    .C(_04103_),
    .Y(_03430_)
  );
  NOR2X1 _10592_ (
    .A(_03969_),
    .B(_04007_),
    .Y(_04104_)
  );
  AOI21X1 _10593_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03970_),
    .C(_04104_),
    .Y(_04105_)
  );
  INVX1 _10594_ (
    .A(_04105_),
    .Y(_04106_)
  );
  NAND2X1 _10595_ (
    .A(_04003_),
    .B(_04106_),
    .Y(_04107_)
  );
  OAI21X1 _10596_ (
    .A(_03747_),
    .B(_04106_),
    .C(_04107_),
    .Y(_03429_)
  );
  NAND2X1 _10597_ (
    .A(_04021_),
    .B(_04106_),
    .Y(_04108_)
  );
  OAI21X1 _10598_ (
    .A(_03748_),
    .B(_04106_),
    .C(_04108_),
    .Y(_03428_)
  );
  NAND2X1 _10599_ (
    .A(_04024_),
    .B(_04106_),
    .Y(_04109_)
  );
  OAI21X1 _10600_ (
    .A(_03749_),
    .B(_04106_),
    .C(_04109_),
    .Y(_03427_)
  );
  NAND2X1 _10601_ (
    .A( execution_unit_0.inst_dext_12_ ),
    .B(_04105_),
    .Y(_04110_)
  );
  OAI21X1 _10602_ (
    .A(_04028_),
    .B(_04105_),
    .C(_04110_),
    .Y(_03426_)
  );
  NAND2X1 _10603_ (
    .A( execution_unit_0.inst_dext_11_ ),
    .B(_04105_),
    .Y(_04111_)
  );
  OAI21X1 _10604_ (
    .A(_04032_),
    .B(_04105_),
    .C(_04111_),
    .Y(_03425_)
  );
  NAND2X1 _10605_ (
    .A( execution_unit_0.inst_dext_10_ ),
    .B(_04105_),
    .Y(_04112_)
  );
  OAI21X1 _10606_ (
    .A(_04038_),
    .B(_04105_),
    .C(_04112_),
    .Y(_03424_)
  );
  NAND2X1 _10607_ (
    .A( execution_unit_0.inst_dext_9_ ),
    .B(_04105_),
    .Y(_04113_)
  );
  OAI21X1 _10608_ (
    .A(_04048_),
    .B(_04105_),
    .C(_04113_),
    .Y(_03423_)
  );
  NAND2X1 _10609_ (
    .A( execution_unit_0.inst_dext_8_ ),
    .B(_04105_),
    .Y(_04114_)
  );
  OAI21X1 _10610_ (
    .A(_04053_),
    .B(_04105_),
    .C(_04114_),
    .Y(_03422_)
  );
  NAND2X1 _10611_ (
    .A( execution_unit_0.inst_dext_7_ ),
    .B(_04105_),
    .Y(_04115_)
  );
  OAI21X1 _10612_ (
    .A(_04058_),
    .B(_04105_),
    .C(_04115_),
    .Y(_03421_)
  );
  NAND2X1 _10613_ (
    .A( execution_unit_0.inst_dext_6_ ),
    .B(_04105_),
    .Y(_04116_)
  );
  OAI21X1 _10614_ (
    .A(_04064_),
    .B(_04105_),
    .C(_04116_),
    .Y(_03420_)
  );
  NAND2X1 _10615_ (
    .A( execution_unit_0.inst_dext_5_ ),
    .B(_04105_),
    .Y(_04117_)
  );
  OAI21X1 _10616_ (
    .A(_04070_),
    .B(_04105_),
    .C(_04117_),
    .Y(_03419_)
  );
  NAND2X1 _10617_ (
    .A(_04078_),
    .B(_04106_),
    .Y(_04118_)
  );
  OAI21X1 _10618_ (
    .A(_03750_),
    .B(_04106_),
    .C(_04118_),
    .Y(_03418_)
  );
  NAND2X1 _10619_ (
    .A( execution_unit_0.inst_dext_3_ ),
    .B(_04105_),
    .Y(_04119_)
  );
  OAI21X1 _10620_ (
    .A(_04082_),
    .B(_04105_),
    .C(_04119_),
    .Y(_03417_)
  );
  NAND2X1 _10621_ (
    .A( execution_unit_0.inst_dext_2_ ),
    .B(_04105_),
    .Y(_04120_)
  );
  OAI21X1 _10622_ (
    .A(_04088_),
    .B(_04105_),
    .C(_04120_),
    .Y(_03416_)
  );
  NAND2X1 _10623_ (
    .A( execution_unit_0.inst_dext_1_ ),
    .B(_04105_),
    .Y(_04121_)
  );
  OAI21X1 _10624_ (
    .A(_04095_),
    .B(_04105_),
    .C(_04121_),
    .Y(_03415_)
  );
  MUX2X1 _10625_ (
    .A( execution_unit_0.inst_dext_0_ ),
    .B( dbg_0.fe_mdb_in_0_ ),
    .S(_04105_),
    .Y(_04122_)
  );
  INVX1 _10626_ (
    .A(_04122_),
    .Y(_03414_)
  );
  OAI21X1 _10627_ (
    .A(_03752_),
    .B(_03911_),
    .C(_03918_),
    .Y(_03413_)
  );
  OAI21X1 _10628_ (
    .A(_03753_),
    .B(_03911_),
    .C(_03965_),
    .Y(_03412_)
  );
  OAI22X1 _10629_ (
    .A(_03754_),
    .B(_03911_),
    .C(_03935_),
    .D(_03909_),
    .Y(_03411_)
  );
  NOR2X1 _10630_ (
    .A(_03766_),
    .B(_03794_),
    .Y(_04123_)
  );
  NAND2X1 _10631_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_04124_)
  );
  NAND3X1 _10632_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03860_),
    .C(_03933_),
    .Y(_04125_)
  );
  NOR2X1 _10633_ (
    .A(_04124_),
    .B(_04125_),
    .Y(_04126_)
  );
  NOR2X1 _10634_ (
    .A(_03859_),
    .B(_04126_),
    .Y(_04127_)
  );
  MUX2X1 _10635_ (
    .A(_03755_),
    .B(_04127_),
    .S(_03910_),
    .Y(_03410_)
  );
  NAND2X1 _10636_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_03910_),
    .Y(_04128_)
  );
  NOR2X1 _10637_ (
    .A(_03766_),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_04129_)
  );
  INVX1 _10638_ (
    .A(_04129_),
    .Y(_04130_)
  );
  NOR2X1 _10639_ (
    .A(_04125_),
    .B(_04130_),
    .Y(_04131_)
  );
  OR2X1 _10640_ (
    .A(_04125_),
    .B(_04130_),
    .Y(_04132_)
  );
  OAI21X1 _10641_ (
    .A(_03910_),
    .B(_04132_),
    .C(_04128_),
    .Y(_03409_)
  );
  NAND2X1 _10642_ (
    .A(_03766_),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_04133_)
  );
  OAI21X1 _10643_ (
    .A(_04125_),
    .B(_04133_),
    .C(_03911_),
    .Y(_04134_)
  );
  OAI21X1 _10644_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_03911_),
    .C(_04134_),
    .Y(_04135_)
  );
  INVX1 _10645_ (
    .A(_04135_),
    .Y(_03408_)
  );
  NAND2X1 _10646_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(_03910_),
    .Y(_04136_)
  );
  OAI21X1 _10647_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03766_),
    .Y(_04137_)
  );
  NOR2X1 _10648_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_04137_),
    .Y(_04138_)
  );
  OR2X1 _10649_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_04137_),
    .Y(_04139_)
  );
  OAI21X1 _10650_ (
    .A(_04125_),
    .B(_04139_),
    .C(_04136_),
    .Y(_03407_)
  );
  NOR2X1 _10651_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03935_),
    .Y(_04140_)
  );
  AOI21X1 _10652_ (
    .A(_04123_),
    .B(_04140_),
    .C(_03910_),
    .Y(_04141_)
  );
  NOR2X1 _10653_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B(_03911_),
    .Y(_04142_)
  );
  NOR2X1 _10654_ (
    .A(_04141_),
    .B(_04142_),
    .Y(_03406_)
  );
  NAND2X1 _10655_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B(_03910_),
    .Y(_04143_)
  );
  NAND3X1 _10656_ (
    .A(_03766_),
    .B( dbg_0.fe_mdb_in_7_ ),
    .C(_04140_),
    .Y(_04144_)
  );
  OAI21X1 _10657_ (
    .A(_03909_),
    .B(_04144_),
    .C(_04143_),
    .Y(_03405_)
  );
  AOI22X1 _10658_ (
    .A( execution_unit_0.alu_0.inst_so_0_ ),
    .B(_03910_),
    .C(_04138_),
    .D(_04140_),
    .Y(_04145_)
  );
  INVX1 _10659_ (
    .A(_04145_),
    .Y(_03404_)
  );
  OAI21X1 _10660_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C( dbg_0.fe_mdb_in_12_ ),
    .Y(_04146_)
  );
  OAI21X1 _10661_ (
    .A(_03757_),
    .B(_03911_),
    .C(_04146_),
    .Y(_03403_)
  );
  MUX2X1 _10662_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .S(_03911_),
    .Y(_04147_)
  );
  INVX1 _10663_ (
    .A(_04147_),
    .Y(_03402_)
  );
  MUX2X1 _10664_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B( frontend_0.inst_jmp_bin_0_ ),
    .S(_03911_),
    .Y(_04148_)
  );
  INVX1 _10665_ (
    .A(_04148_),
    .Y(_03401_)
  );
  NAND2X1 _10666_ (
    .A( execution_unit_0.inst_mov ),
    .B(_03910_),
    .Y(_04149_)
  );
  NAND3X1 _10667_ (
    .A(_03756_),
    .B( dbg_0.fe_mdb_in_14_ ),
    .C(_03791_),
    .Y(_04150_)
  );
  OR2X1 _10668_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_04150_),
    .Y(_04151_)
  );
  OAI21X1 _10669_ (
    .A(_03918_),
    .B(_04151_),
    .C(_04149_),
    .Y(_03400_)
  );
  OAI21X1 _10670_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03759_),
    .Y(_04152_)
  );
  OAI21X1 _10671_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03911_),
    .C(_04152_),
    .Y(_04153_)
  );
  INVX1 _10672_ (
    .A(_04153_),
    .Y(_03399_)
  );
  MUX2X1 _10673_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .S(_03911_),
    .Y(_04154_)
  );
  INVX1 _10674_ (
    .A(_04154_),
    .Y(_03398_)
  );
  OAI21X1 _10675_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03762_),
    .Y(_04155_)
  );
  OAI21X1 _10676_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B(_03911_),
    .C(_04155_),
    .Y(_04156_)
  );
  INVX1 _10677_ (
    .A(_04156_),
    .Y(_03397_)
  );
  OAI21X1 _10678_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03751_),
    .Y(_04157_)
  );
  OAI21X1 _10679_ (
    .A( frontend_0.inst_dest_bin_0_ ),
    .B(_03911_),
    .C(_04157_),
    .Y(_04158_)
  );
  INVX1 _10680_ (
    .A(_04158_),
    .Y(_03396_)
  );
  OAI21X1 _10681_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_03764_),
    .Y(_04159_)
  );
  OAI21X1 _10682_ (
    .A( frontend_0.inst_src_bin_1_ ),
    .B(_03911_),
    .C(_04159_),
    .Y(_04160_)
  );
  INVX1 _10683_ (
    .A(_04160_),
    .Y(_03395_)
  );
  OAI21X1 _10684_ (
    .A( frontend_0.inst_src_bin_0_ ),
    .B(_03911_),
    .C(_04137_),
    .Y(_04161_)
  );
  INVX1 _10685_ (
    .A(_04161_),
    .Y(_03394_)
  );
  OAI21X1 _10686_ (
    .A(_03768_),
    .B(_03911_),
    .C(_03963_),
    .Y(_03393_)
  );
  NAND2X1 _10687_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B(_03910_),
    .Y(_04162_)
  );
  NAND3X1 _10688_ (
    .A(_03792_),
    .B( dbg_0.fe_mdb_in_4_ ),
    .C(_03932_),
    .Y(_04163_)
  );
  OR2X1 _10689_ (
    .A(_03910_),
    .B(_04163_),
    .Y(_04164_)
  );
  OAI21X1 _10690_ (
    .A(_03959_),
    .B(_04164_),
    .C(_04162_),
    .Y(_03392_)
  );
  NAND2X1 _10691_ (
    .A(_03946_),
    .B(_03957_),
    .Y(_04165_)
  );
  NOR3X1 _10692_ (
    .A(_03947_),
    .B(_03958_),
    .C(_04015_),
    .Y(_04166_)
  );
  NAND3X1 _10693_ (
    .A(_03946_),
    .B(_03957_),
    .C(_04014_),
    .Y(_04167_)
  );
  OAI21X1 _10694_ (
    .A(_03859_),
    .B( dbg_0.decode_noirq ),
    .C(_04167_),
    .Y(_04168_)
  );
  OAI21X1 _10695_ (
    .A( execution_unit_0.inst_as_5_ ),
    .B(_03911_),
    .C(_04168_),
    .Y(_04169_)
  );
  INVX1 _10696_ (
    .A(_04169_),
    .Y(_03391_)
  );
  OAI22X1 _10697_ (
    .A(_03769_),
    .B(_03911_),
    .C(_04164_),
    .D(_04165_),
    .Y(_03390_)
  );
  NAND2X1 _10698_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B(_03910_),
    .Y(_04170_)
  );
  NAND2X1 _10699_ (
    .A(_03949_),
    .B(_03958_),
    .Y(_04171_)
  );
  NOR3X1 _10700_ (
    .A(_03948_),
    .B(_03957_),
    .C(_04015_),
    .Y(_04172_)
  );
  NAND3X1 _10701_ (
    .A(_03949_),
    .B(_03958_),
    .C(_04014_),
    .Y(_04173_)
  );
  OAI21X1 _10702_ (
    .A(_03910_),
    .B(_04173_),
    .C(_04170_),
    .Y(_03389_)
  );
  OAI21X1 _10703_ (
    .A(_03948_),
    .B(_04091_),
    .C(_03911_),
    .Y(_04174_)
  );
  OAI21X1 _10704_ (
    .A( execution_unit_0.inst_as_2_ ),
    .B(_03911_),
    .C(_04174_),
    .Y(_04175_)
  );
  INVX1 _10705_ (
    .A(_04175_),
    .Y(_03388_)
  );
  NAND2X1 _10706_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B(_03910_),
    .Y(_04176_)
  );
  OAI21X1 _10707_ (
    .A(_04164_),
    .B(_04171_),
    .C(_04176_),
    .Y(_03387_)
  );
  NAND2X1 _10708_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B(_03910_),
    .Y(_04177_)
  );
  NAND3X1 _10709_ (
    .A(_03956_),
    .B(_03960_),
    .C(_04013_),
    .Y(_04178_)
  );
  OAI21X1 _10710_ (
    .A(_03910_),
    .B(_04178_),
    .C(_04177_),
    .Y(_03386_)
  );
  NAND2X1 _10711_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_03910_),
    .Y(_04179_)
  );
  NAND3X1 _10712_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03854_),
    .C(_03932_),
    .Y(_04180_)
  );
  OAI21X1 _10713_ (
    .A(_03915_),
    .B(_04180_),
    .C(_04179_),
    .Y(_03385_)
  );
  AOI21X1 _10714_ (
    .A(_03948_),
    .B(_03954_),
    .C(_04163_),
    .Y(_04181_)
  );
  NOR2X1 _10715_ (
    .A(_04166_),
    .B(_04181_),
    .Y(_04182_)
  );
  OAI21X1 _10716_ (
    .A(_03925_),
    .B(_04182_),
    .C(_03911_),
    .Y(_04183_)
  );
  OAI21X1 _10717_ (
    .A( frontend_0.inst_sz_1_ ),
    .B(_03911_),
    .C(_04183_),
    .Y(_04184_)
  );
  INVX1 _10718_ (
    .A(_04184_),
    .Y(_03384_)
  );
  AND2X1 _10719_ (
    .A(_03925_),
    .B(_04182_),
    .Y(_04185_)
  );
  NAND2X1 _10720_ (
    .A( frontend_0.inst_sz_0_ ),
    .B(_03910_),
    .Y(_04186_)
  );
  OAI21X1 _10721_ (
    .A(_04183_),
    .B(_04185_),
    .C(_04186_),
    .Y(_03383_)
  );
  AOI21X1 _10722_ (
    .A(_03923_),
    .B(_03930_),
    .C(_03824_),
    .Y(_04187_)
  );
  AOI21X1 _10723_ (
    .A(_03911_),
    .B(_04131_),
    .C(_03964_),
    .Y(_04188_)
  );
  NAND2X1 _10724_ (
    .A(_04187_),
    .B(_04188_),
    .Y(_03382_)
  );
  OR2X1 _10725_ (
    .A(_03825_),
    .B(_03906_),
    .Y(_04189_)
  );
  OAI21X1 _10726_ (
    .A(_03772_),
    .B(_03827_),
    .C(_04189_),
    .Y(_03381_)
  );
  NOR2X1 _10727_ (
    .A(_03826_),
    .B(_03831_),
    .Y(_04190_)
  );
  NAND2X1 _10728_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B(_04190_),
    .Y(_04191_)
  );
  OAI21X1 _10729_ (
    .A(_03830_),
    .B(_03831_),
    .C( frontend_0.exec_src_wr ),
    .Y(_04192_)
  );
  OAI21X1 _10730_ (
    .A(_03827_),
    .B(_04192_),
    .C(_04191_),
    .Y(_03380_)
  );
  OAI21X1 _10731_ (
    .A( frontend_0.exec_dext_rdy ),
    .B(_04106_),
    .C(_04189_),
    .Y(_04193_)
  );
  INVX1 _10732_ (
    .A(_04193_),
    .Y(_03379_)
  );
  NAND2X1 _10733_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_03910_),
    .Y(_04194_)
  );
  AND2X1 _10734_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03860_),
    .Y(_04195_)
  );
  NAND2X1 _10735_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03860_),
    .Y(_04196_)
  );
  NAND2X1 _10736_ (
    .A(_03790_),
    .B(_04195_),
    .Y(_04197_)
  );
  OAI21X1 _10737_ (
    .A(_04146_),
    .B(_04197_),
    .C(_04194_),
    .Y(_03378_)
  );
  NAND3X1 _10738_ (
    .A(_03794_),
    .B(_03911_),
    .C(_04140_),
    .Y(_04198_)
  );
  OAI21X1 _10739_ (
    .A(_03774_),
    .B(_03911_),
    .C(_04198_),
    .Y(_03377_)
  );
  NAND2X1 _10740_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B( dbg_0.fe_mdb_in_14_ ),
    .Y(_04199_)
  );
  NOR2X1 _10741_ (
    .A(_03756_),
    .B(_03791_),
    .Y(_04200_)
  );
  NOR2X1 _10742_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03859_),
    .Y(_03455_)
  );
  NAND3X1 _10743_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_04200_),
    .C(_03455_),
    .Y(_03456_)
  );
  OR2X1 _10744_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_04197_),
    .Y(_03457_)
  );
  OAI21X1 _10745_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_04197_),
    .C(_03456_),
    .Y(_03458_)
  );
  NOR2X1 _10746_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B(_03791_),
    .Y(_03459_)
  );
  AND2X1 _10747_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03459_),
    .Y(_03460_)
  );
  NAND2X1 _10748_ (
    .A(_03455_),
    .B(_03460_),
    .Y(_03461_)
  );
  NOR2X1 _10749_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_04199_),
    .Y(_03462_)
  );
  OAI21X1 _10750_ (
    .A(_03460_),
    .B(_03462_),
    .C(_03455_),
    .Y(_03463_)
  );
  INVX1 _10751_ (
    .A(_03463_),
    .Y(_03464_)
  );
  OAI21X1 _10752_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03794_),
    .C(_04140_),
    .Y(_03465_)
  );
  NAND2X1 _10753_ (
    .A(_04195_),
    .B(_03460_),
    .Y(_03466_)
  );
  AOI21X1 _10754_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_04195_),
    .C(_03910_),
    .Y(_03467_)
  );
  OAI21X1 _10755_ (
    .A(_03458_),
    .B(_03464_),
    .C(_03911_),
    .Y(_03468_)
  );
  NAND3X1 _10756_ (
    .A(_03465_),
    .B(_03467_),
    .C(_03468_),
    .Y(_03469_)
  );
  OAI21X1 _10757_ (
    .A( execution_unit_0.alu_0.inst_alu_9_ ),
    .B(_03911_),
    .C(_03469_),
    .Y(_03470_)
  );
  INVX1 _10758_ (
    .A(_03470_),
    .Y(_03376_)
  );
  NAND2X1 _10759_ (
    .A(_04195_),
    .B(_04200_),
    .Y(_03471_)
  );
  NOR2X1 _10760_ (
    .A( execution_unit_0.alu_0.inst_alu_8_ ),
    .B(_03911_),
    .Y(_03472_)
  );
  AOI21X1 _10761_ (
    .A(_04141_),
    .B(_03471_),
    .C(_03472_),
    .Y(_03375_)
  );
  NAND3X1 _10762_ (
    .A(_03790_),
    .B(_04195_),
    .C(_03459_),
    .Y(_03473_)
  );
  NAND2X1 _10763_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_03910_),
    .Y(_03474_)
  );
  OAI21X1 _10764_ (
    .A(_03909_),
    .B(_03473_),
    .C(_03474_),
    .Y(_03374_)
  );
  NAND2X1 _10765_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_03910_),
    .Y(_03475_)
  );
  OAI21X1 _10766_ (
    .A(_03909_),
    .B(_03466_),
    .C(_03475_),
    .Y(_03373_)
  );
  NAND2X1 _10767_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_03910_),
    .Y(_03476_)
  );
  NAND2X1 _10768_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03462_),
    .Y(_03477_)
  );
  OAI21X1 _10769_ (
    .A(_03915_),
    .B(_03477_),
    .C(_03476_),
    .Y(_03372_)
  );
  OAI21X1 _10770_ (
    .A(_04150_),
    .B(_04196_),
    .C(_03911_),
    .Y(_03478_)
  );
  INVX1 _10771_ (
    .A(_03478_),
    .Y(_03479_)
  );
  NOR2X1 _10772_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_03911_),
    .Y(_03480_)
  );
  AOI21X1 _10773_ (
    .A(_03471_),
    .B(_03479_),
    .C(_03480_),
    .Y(_03371_)
  );
  NAND2X1 _10774_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_03910_),
    .Y(_03481_)
  );
  NAND3X1 _10775_ (
    .A(_04188_),
    .B(_03468_),
    .C(_03481_),
    .Y(_03370_)
  );
  NAND3X1 _10776_ (
    .A(_03456_),
    .B(_03461_),
    .C(_03473_),
    .Y(_03482_)
  );
  MUX2X1 _10777_ (
    .A( execution_unit_0.alu_0.inst_alu_2_ ),
    .B(_03482_),
    .S(_03910_),
    .Y(_03483_)
  );
  INVX1 _10778_ (
    .A(_03483_),
    .Y(_03369_)
  );
  NAND2X1 _10779_ (
    .A( execution_unit_0.alu_0.inst_alu_1_ ),
    .B(_03910_),
    .Y(_03484_)
  );
  OAI21X1 _10780_ (
    .A(_03909_),
    .B(_03457_),
    .C(_03484_),
    .Y(_03368_)
  );
  OAI22X1 _10781_ (
    .A( execution_unit_0.alu_0.inst_alu_0_ ),
    .B(_03911_),
    .C(_03458_),
    .D(_03478_),
    .Y(_03485_)
  );
  INVX1 _10782_ (
    .A(_03485_),
    .Y(_03367_)
  );
  AOI21X1 _10783_ (
    .A(_03949_),
    .B(_04090_),
    .C(_04131_),
    .Y(_03486_)
  );
  OAI21X1 _10784_ (
    .A(_03948_),
    .B(_04091_),
    .C(_04132_),
    .Y(_03487_)
  );
  NOR3X1 _10785_ (
    .A(_04166_),
    .B(_04172_),
    .C(_03487_),
    .Y(_03488_)
  );
  NAND3X1 _10786_ (
    .A(_04167_),
    .B(_04173_),
    .C(_03486_),
    .Y(_03489_)
  );
  NOR2X1 _10787_ (
    .A( clock_module_0.UNUSED_cpuoff ),
    .B(_03855_),
    .Y(_03490_)
  );
  OAI21X1 _10788_ (
    .A(_03778_),
    .B(_03818_),
    .C(_03490_),
    .Y(_03491_)
  );
  INVX1 _10789_ (
    .A(_03491_),
    .Y(_03492_)
  );
  NOR2X1 _10790_ (
    .A(_04181_),
    .B(_03491_),
    .Y(_03493_)
  );
  OAI21X1 _10791_ (
    .A(_03955_),
    .B(_04163_),
    .C(_03492_),
    .Y(_03494_)
  );
  OAI21X1 _10792_ (
    .A(_03924_),
    .B(_03489_),
    .C(_03493_),
    .Y(_03495_)
  );
  NOR2X1 _10793_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_04127_),
    .Y(_03496_)
  );
  OAI21X1 _10794_ (
    .A(_03859_),
    .B(_04126_),
    .C(_03786_),
    .Y(_03497_)
  );
  NAND2X1 _10795_ (
    .A(_03772_),
    .B(_03834_),
    .Y(_03498_)
  );
  NOR2X1 _10796_ (
    .A( frontend_0.exec_jmp ),
    .B(_03498_),
    .Y(_03499_)
  );
  OAI21X1 _10797_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_03822_),
    .C(_03833_),
    .Y(_03500_)
  );
  NOR2X1 _10798_ (
    .A(_03827_),
    .B(_03500_),
    .Y(_03501_)
  );
  AOI21X1 _10799_ (
    .A(_03771_),
    .B(_03827_),
    .C(_03500_),
    .Y(_03502_)
  );
  OAI21X1 _10800_ (
    .A( frontend_0.exec_jmp ),
    .B(_03498_),
    .C(_03502_),
    .Y(_03503_)
  );
  AND2X1 _10801_ (
    .A(_03497_),
    .B(_03503_),
    .Y(_03504_)
  );
  NOR2X1 _10802_ (
    .A(_03821_),
    .B(_03825_),
    .Y(_03505_)
  );
  OAI21X1 _10803_ (
    .A( frontend_0.exec_dext_rdy ),
    .B(_04106_),
    .C(_03505_),
    .Y(_03506_)
  );
  OR2X1 _10804_ (
    .A(_03831_),
    .B(_03906_),
    .Y(_03507_)
  );
  OR2X1 _10805_ (
    .A( execution_unit_0.inst_ad_6_ ),
    .B( execution_unit_0.UNUSED_inst_ad_symb ),
    .Y(_03508_)
  );
  NOR2X1 _10806_ (
    .A( execution_unit_0.UNUSED_inst_ad_idx ),
    .B(_03508_),
    .Y(_03509_)
  );
  AND2X1 _10807_ (
    .A(_04190_),
    .B(_03509_),
    .Y(_03510_)
  );
  NAND2X1 _10808_ (
    .A(_03788_),
    .B(_03789_),
    .Y(_03511_)
  );
  OAI21X1 _10809_ (
    .A(_03821_),
    .B(_03831_),
    .C(_04189_),
    .Y(_03512_)
  );
  INVX1 _10810_ (
    .A(_03512_),
    .Y(_03513_)
  );
  OAI21X1 _10811_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03511_),
    .C(_03513_),
    .Y(_03514_)
  );
  NOR2X1 _10812_ (
    .A(_03510_),
    .B(_03514_),
    .Y(_03515_)
  );
  OAI21X1 _10813_ (
    .A(_04009_),
    .B(_03507_),
    .C(_03515_),
    .Y(_03516_)
  );
  AOI21X1 _10814_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03499_),
    .C(_03516_),
    .Y(_03517_)
  );
  NAND2X1 _10815_ (
    .A(_03506_),
    .B(_03517_),
    .Y(_03518_)
  );
  AOI21X1 _10816_ (
    .A(_03495_),
    .B(_03504_),
    .C(_03518_),
    .Y(_03519_)
  );
  INVX1 _10817_ (
    .A(_03519_),
    .Y( frontend_0.e_state_nxt_0_ )
  );
  OAI21X1 _10818_ (
    .A( frontend_0.exec_dst_wr ),
    .B(_03835_),
    .C(_03501_),
    .Y(_03520_)
  );
  OAI21X1 _10819_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_04127_),
    .C(_03520_),
    .Y(_03521_)
  );
  AOI21X1 _10820_ (
    .A(_03488_),
    .B(_03493_),
    .C(_03521_),
    .Y(_03522_)
  );
  OAI21X1 _10821_ (
    .A(_03830_),
    .B(_03511_),
    .C(_03507_),
    .Y(_03523_)
  );
  AOI21X1 _10822_ (
    .A( frontend_0.exec_jmp ),
    .B(_03827_),
    .C(_03523_),
    .Y(_03524_)
  );
  NOR2X1 _10823_ (
    .A( frontend_0.exec_jmp ),
    .B( frontend_0.exec_src_wr ),
    .Y(_03525_)
  );
  OAI21X1 _10824_ (
    .A(_03498_),
    .B(_03525_),
    .C(_03524_),
    .Y(_03526_)
  );
  NOR2X1 _10825_ (
    .A(_03522_),
    .B(_03526_),
    .Y(_03527_)
  );
  INVX1 _10826_ (
    .A(_03527_),
    .Y( frontend_0.e_state_nxt_2_ )
  );
  OAI21X1 _10827_ (
    .A(_04181_),
    .B(_03489_),
    .C(_03492_),
    .Y(_03528_)
  );
  OAI21X1 _10828_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03835_),
    .C(_03501_),
    .Y(_03529_)
  );
  AND2X1 _10829_ (
    .A(_03497_),
    .B(_03529_),
    .Y(_03530_)
  );
  OAI22X1 _10830_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_03825_),
    .C(_03831_),
    .D( execution_unit_0.e_state_0_ ),
    .Y(_03531_)
  );
  AOI21X1 _10831_ (
    .A( frontend_0.exec_jmp ),
    .B(_03827_),
    .C(_03834_),
    .Y(_03532_)
  );
  AOI21X1 _10832_ (
    .A(_03771_),
    .B(_03772_),
    .C(_03532_),
    .Y(_03533_)
  );
  OR2X1 _10833_ (
    .A(_03531_),
    .B(_03533_),
    .Y(_03534_)
  );
  AOI21X1 _10834_ (
    .A(_03528_),
    .B(_03530_),
    .C(_03534_),
    .Y(_03535_)
  );
  INVX1 _10835_ (
    .A(_03535_),
    .Y( frontend_0.e_state_nxt_3_ )
  );
  NAND2X1 _10836_ (
    .A(_03795_),
    .B(_03916_),
    .Y(_03536_)
  );
  NOR2X1 _10837_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03971_),
    .Y(_03537_)
  );
  NAND2X1 _10838_ (
    .A(_03778_),
    .B(_03970_),
    .Y(_03538_)
  );
  OAI21X1 _10839_ (
    .A(_03854_),
    .B(_03907_),
    .C(_03838_),
    .Y(_03539_)
  );
  OAI21X1 _10840_ (
    .A( clock_module_0.UNUSED_cpuoff ),
    .B(_03855_),
    .C(_03539_),
    .Y(_03540_)
  );
  NOR2X1 _10841_ (
    .A(_03905_),
    .B(_03540_),
    .Y(_03541_)
  );
  NOR2X1 _10842_ (
    .A(_03820_),
    .B(_03490_),
    .Y(_03542_)
  );
  AOI22X1 _10843_ (
    .A(_03860_),
    .B(_03541_),
    .C(_03542_),
    .D(_03858_),
    .Y(_03543_)
  );
  AND2X1 _10844_ (
    .A(_03538_),
    .B(_03543_),
    .Y(_03544_)
  );
  OAI21X1 _10845_ (
    .A(_04185_),
    .B(_03536_),
    .C(_03544_),
    .Y( frontend_0.i_state_nxt_0_ )
  );
  OAI21X1 _10846_ (
    .A(_03969_),
    .B(_03974_),
    .C(_03543_),
    .Y( frontend_0.i_state_nxt_2_ )
  );
  AOI22X1 _10847_ (
    .A(_03819_),
    .B(_03490_),
    .C(_03540_),
    .D(_03904_),
    .Y(_03545_)
  );
  NOR2X1 _10848_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03818_),
    .Y(_03546_)
  );
  NAND2X1 _10849_ (
    .A(_03778_),
    .B(_03817_),
    .Y(_03547_)
  );
  NAND3X1 _10850_ (
    .A(_03972_),
    .B(_03975_),
    .C(_03547_),
    .Y(_03548_)
  );
  INVX1 _10851_ (
    .A(_03548_),
    .Y(_03549_)
  );
  OAI21X1 _10852_ (
    .A(_03859_),
    .B(_03545_),
    .C(_03549_),
    .Y( frontend_0.i_state_nxt_1_ )
  );
  OAI21X1 _10853_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_04125_),
    .C(_03925_),
    .Y(_03550_)
  );
  AOI21X1 _10854_ (
    .A(_03488_),
    .B(_03550_),
    .C(_03494_),
    .Y(_03551_)
  );
  NOR2X1 _10855_ (
    .A(_03496_),
    .B(_03551_),
    .Y(_03552_)
  );
  AOI21X1 _10856_ (
    .A(_03773_),
    .B(_03552_),
    .C( frontend_0.exec_jmp ),
    .Y(_03553_)
  );
  OAI21X1 _10857_ (
    .A( frontend_0.exec_dst_wr ),
    .B(_03553_),
    .C(_03834_),
    .Y(_03554_)
  );
  OR2X1 _10858_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_03555_)
  );
  OR2X1 _10859_ (
    .A( execution_unit_0.UNUSED_inst_ad_idx ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_03556_)
  );
  NOR2X1 _10860_ (
    .A(_03555_),
    .B(_03556_),
    .Y(_03557_)
  );
  OAI22X1 _10861_ (
    .A(_03787_),
    .B(_03822_),
    .C(_03511_),
    .D(_03821_),
    .Y(_03558_)
  );
  NOR2X1 _10862_ (
    .A(_03512_),
    .B(_03558_),
    .Y(_03559_)
  );
  OAI21X1 _10863_ (
    .A(_04008_),
    .B(_03507_),
    .C(_03559_),
    .Y(_03560_)
  );
  AOI21X1 _10864_ (
    .A(_03510_),
    .B(_03557_),
    .C(_03560_),
    .Y(_03561_)
  );
  OAI21X1 _10865_ (
    .A(_03502_),
    .B(_03552_),
    .C(_03561_),
    .Y(_03562_)
  );
  INVX1 _10866_ (
    .A(_03562_),
    .Y(_03563_)
  );
  NAND2X1 _10867_ (
    .A(_03554_),
    .B(_03563_),
    .Y( frontend_0.e_state_nxt_1_ )
  );
  OAI21X1 _10868_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03971_),
    .C(_03795_),
    .Y(_03564_)
  );
  AOI21X1 _10869_ (
    .A(_03751_),
    .B(_03546_),
    .C(_03564_),
    .Y(_03565_)
  );
  OAI21X1 _10870_ (
    .A( dbg_0.UNUSED_pc_0_ ),
    .B(_03546_),
    .C(_03565_),
    .Y(_03566_)
  );
  OAI21X1 _10871_ (
    .A(_03795_),
    .B(_03796_),
    .C(_03566_),
    .Y( execution_unit_0.pc_nxt_0_ )
  );
  NOR2X1 _10872_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_03567_)
  );
  NOR2X1 _10873_ (
    .A(_03905_),
    .B(_03908_),
    .Y(_03568_)
  );
  OR2X1 _10874_ (
    .A(_03905_),
    .B(_03908_),
    .Y(_03569_)
  );
  NOR3X1 _10875_ (
    .A(_03519_),
    .B(_03527_),
    .C(_03535_),
    .Y(_03570_)
  );
  NAND3X1 _10876_ (
    .A( frontend_0.e_state_nxt_0_ ),
    .B( frontend_0.e_state_nxt_2_ ),
    .C( frontend_0.e_state_nxt_3_ ),
    .Y(_03571_)
  );
  OAI21X1 _10877_ (
    .A(_03568_),
    .B(_03570_),
    .C(_03797_),
    .Y(_03572_)
  );
  NOR3X1 _10878_ (
    .A(_03797_),
    .B(_03568_),
    .C(_03570_),
    .Y(_03573_)
  );
  NAND3X1 _10879_ (
    .A( dbg_0.UNUSED_pc_1_ ),
    .B(_03569_),
    .C(_03571_),
    .Y(_03574_)
  );
  NAND2X1 _10880_ (
    .A(_03572_),
    .B(_03574_),
    .Y(_03575_)
  );
  OAI21X1 _10881_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B(_03547_),
    .C(_03538_),
    .Y(_03576_)
  );
  AOI21X1 _10882_ (
    .A(_03547_),
    .B(_03575_),
    .C(_03576_),
    .Y(_03577_)
  );
  AOI21X1 _10883_ (
    .A( frontend_0.irq_addr_1_ ),
    .B(_03537_),
    .C(_03577_),
    .Y(_03578_)
  );
  AOI21X1 _10884_ (
    .A(_03795_),
    .B(_03578_),
    .C(_03567_),
    .Y( execution_unit_0.pc_nxt_1_ )
  );
  NOR2X1 _10885_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_03579_)
  );
  XNOR2X1 _10886_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .B(_03573_),
    .Y(_03580_)
  );
  AOI21X1 _10887_ (
    .A(_03547_),
    .B(_03580_),
    .C(_03537_),
    .Y(_03581_)
  );
  OAI21X1 _10888_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_03547_),
    .C(_03581_),
    .Y(_03582_)
  );
  AOI21X1 _10889_ (
    .A( frontend_0.irq_addr_2_ ),
    .B(_03537_),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03583_)
  );
  AOI21X1 _10890_ (
    .A(_03582_),
    .B(_03583_),
    .C(_03579_),
    .Y( execution_unit_0.pc_nxt_2_ )
  );
  NOR2X1 _10891_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_03584_)
  );
  AOI21X1 _10892_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .B(_03573_),
    .C( dbg_0.UNUSED_pc_3_ ),
    .Y(_03585_)
  );
  NOR3X1 _10893_ (
    .A(_03798_),
    .B(_03799_),
    .C(_03574_),
    .Y(_03586_)
  );
  NAND3X1 _10894_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .B( dbg_0.UNUSED_pc_3_ ),
    .C(_03573_),
    .Y(_03587_)
  );
  OAI21X1 _10895_ (
    .A(_03585_),
    .B(_03586_),
    .C(_03547_),
    .Y(_03588_)
  );
  AOI21X1 _10896_ (
    .A(_03759_),
    .B(_03546_),
    .C(_03537_),
    .Y(_03589_)
  );
  OAI21X1 _10897_ (
    .A(_03743_),
    .B(_03538_),
    .C(_03795_),
    .Y(_03590_)
  );
  AOI21X1 _10898_ (
    .A(_03588_),
    .B(_03589_),
    .C(_03590_),
    .Y(_03591_)
  );
  NOR2X1 _10899_ (
    .A(_03584_),
    .B(_03591_),
    .Y( execution_unit_0.pc_nxt_3_ )
  );
  NOR2X1 _10900_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_03592_)
  );
  XNOR2X1 _10901_ (
    .A(_03800_),
    .B(_03586_),
    .Y(_03593_)
  );
  AOI21X1 _10902_ (
    .A(_03793_),
    .B(_03546_),
    .C(_03537_),
    .Y(_03594_)
  );
  OAI21X1 _10903_ (
    .A(_03546_),
    .B(_03593_),
    .C(_03594_),
    .Y(_03595_)
  );
  NAND2X1 _10904_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03537_),
    .Y(_03596_)
  );
  AOI21X1 _10905_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03537_),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03597_)
  );
  AOI21X1 _10906_ (
    .A(_03595_),
    .B(_03597_),
    .C(_03592_),
    .Y( execution_unit_0.pc_nxt_4_ )
  );
  NOR3X1 _10907_ (
    .A(_03800_),
    .B(_03801_),
    .C(_03587_),
    .Y(_03598_)
  );
  NAND3X1 _10908_ (
    .A( dbg_0.UNUSED_pc_4_ ),
    .B( dbg_0.UNUSED_pc_5_ ),
    .C(_03586_),
    .Y(_03599_)
  );
  OAI21X1 _10909_ (
    .A(_03800_),
    .B(_03587_),
    .C(_03801_),
    .Y(_03600_)
  );
  OAI21X1 _10910_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03818_),
    .C(_03600_),
    .Y(_03601_)
  );
  AOI21X1 _10911_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03602_)
  );
  OAI21X1 _10912_ (
    .A(_03598_),
    .B(_03601_),
    .C(_03602_),
    .Y(_03603_)
  );
  OAI21X1 _10913_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_5_ ),
    .C(_03603_),
    .Y(_03604_)
  );
  INVX1 _10914_ (
    .A(_03604_),
    .Y( execution_unit_0.pc_nxt_5_ )
  );
  NOR2X1 _10915_ (
    .A(_03802_),
    .B(_03599_),
    .Y(_03605_)
  );
  OAI21X1 _10916_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B(_03598_),
    .C(_03547_),
    .Y(_03606_)
  );
  AOI21X1 _10917_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03607_)
  );
  OAI21X1 _10918_ (
    .A(_03605_),
    .B(_03606_),
    .C(_03607_),
    .Y(_03608_)
  );
  OAI21X1 _10919_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .C(_03608_),
    .Y(_03609_)
  );
  INVX1 _10920_ (
    .A(_03609_),
    .Y( execution_unit_0.pc_nxt_6_ )
  );
  NOR3X1 _10921_ (
    .A(_03802_),
    .B(_03804_),
    .C(_03599_),
    .Y(_03610_)
  );
  NAND3X1 _10922_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B( dbg_0.UNUSED_pc_7_ ),
    .C(_03598_),
    .Y(_03611_)
  );
  OAI21X1 _10923_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .B(_03605_),
    .C(_03547_),
    .Y(_03612_)
  );
  AOI21X1 _10924_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03613_)
  );
  OAI21X1 _10925_ (
    .A(_03610_),
    .B(_03612_),
    .C(_03613_),
    .Y(_03614_)
  );
  OAI21X1 _10926_ (
    .A(_03795_),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .C(_03614_),
    .Y(_03615_)
  );
  INVX1 _10927_ (
    .A(_03615_),
    .Y( execution_unit_0.pc_nxt_7_ )
  );
  XNOR2X1 _10928_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .B(_03610_),
    .Y(_03616_)
  );
  AOI21X1 _10929_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03617_)
  );
  OAI21X1 _10930_ (
    .A(_03546_),
    .B(_03616_),
    .C(_03617_),
    .Y(_03618_)
  );
  OAI21X1 _10931_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_8_ ),
    .C(_03618_),
    .Y(_03619_)
  );
  INVX1 _10932_ (
    .A(_03619_),
    .Y( execution_unit_0.pc_nxt_8_ )
  );
  NOR3X1 _10933_ (
    .A(_03805_),
    .B(_03806_),
    .C(_03611_),
    .Y(_03620_)
  );
  NAND3X1 _10934_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .B( dbg_0.UNUSED_pc_9_ ),
    .C(_03610_),
    .Y(_03621_)
  );
  OAI21X1 _10935_ (
    .A(_03805_),
    .B(_03611_),
    .C(_03806_),
    .Y(_03622_)
  );
  OAI21X1 _10936_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03818_),
    .C(_03622_),
    .Y(_03623_)
  );
  AOI21X1 _10937_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03624_)
  );
  OAI21X1 _10938_ (
    .A(_03620_),
    .B(_03623_),
    .C(_03624_),
    .Y(_03625_)
  );
  OAI21X1 _10939_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_9_ ),
    .C(_03625_),
    .Y(_03626_)
  );
  INVX1 _10940_ (
    .A(_03626_),
    .Y( execution_unit_0.pc_nxt_9_ )
  );
  NOR2X1 _10941_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_10_ ),
    .Y(_03627_)
  );
  AOI21X1 _10942_ (
    .A(_03807_),
    .B(_03621_),
    .C(_03546_),
    .Y(_03628_)
  );
  OAI21X1 _10943_ (
    .A(_03807_),
    .B(_03621_),
    .C(_03628_),
    .Y(_03629_)
  );
  AOI21X1 _10944_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03630_)
  );
  AOI21X1 _10945_ (
    .A(_03629_),
    .B(_03630_),
    .C(_03627_),
    .Y( execution_unit_0.pc_nxt_10_ )
  );
  NOR2X1 _10946_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_11_ ),
    .Y(_03631_)
  );
  NOR3X1 _10947_ (
    .A(_03807_),
    .B(_03808_),
    .C(_03621_),
    .Y(_03632_)
  );
  NAND3X1 _10948_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .B( dbg_0.UNUSED_pc_11_ ),
    .C(_03620_),
    .Y(_03633_)
  );
  OAI21X1 _10949_ (
    .A(_03807_),
    .B(_03621_),
    .C(_03808_),
    .Y(_03634_)
  );
  NAND3X1 _10950_ (
    .A(_03547_),
    .B(_03633_),
    .C(_03634_),
    .Y(_03635_)
  );
  AOI21X1 _10951_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03636_)
  );
  AOI21X1 _10952_ (
    .A(_03635_),
    .B(_03636_),
    .C(_03631_),
    .Y( execution_unit_0.pc_nxt_11_ )
  );
  XNOR2X1 _10953_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .B(_03632_),
    .Y(_03637_)
  );
  AOI21X1 _10954_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03638_)
  );
  OAI21X1 _10955_ (
    .A(_03546_),
    .B(_03637_),
    .C(_03638_),
    .Y(_03639_)
  );
  OAI21X1 _10956_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_12_ ),
    .C(_03639_),
    .Y(_03640_)
  );
  INVX1 _10957_ (
    .A(_03640_),
    .Y( execution_unit_0.pc_nxt_12_ )
  );
  NOR2X1 _10958_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_13_ ),
    .Y(_03641_)
  );
  NOR3X1 _10959_ (
    .A(_03809_),
    .B(_03810_),
    .C(_03633_),
    .Y(_03642_)
  );
  NAND3X1 _10960_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .B( dbg_0.UNUSED_pc_13_ ),
    .C(_03632_),
    .Y(_03643_)
  );
  OAI21X1 _10961_ (
    .A(_03809_),
    .B(_03633_),
    .C(_03810_),
    .Y(_03644_)
  );
  NAND3X1 _10962_ (
    .A(_03547_),
    .B(_03643_),
    .C(_03644_),
    .Y(_03645_)
  );
  AOI21X1 _10963_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03646_)
  );
  AOI21X1 _10964_ (
    .A(_03645_),
    .B(_03646_),
    .C(_03641_),
    .Y( execution_unit_0.pc_nxt_13_ )
  );
  NOR2X1 _10965_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_14_ ),
    .Y(_03647_)
  );
  AOI21X1 _10966_ (
    .A(_03811_),
    .B(_03643_),
    .C(_03546_),
    .Y(_03648_)
  );
  OAI21X1 _10967_ (
    .A(_03811_),
    .B(_03643_),
    .C(_03648_),
    .Y(_03649_)
  );
  AOI21X1 _10968_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03650_)
  );
  AOI21X1 _10969_ (
    .A(_03649_),
    .B(_03650_),
    .C(_03647_),
    .Y( execution_unit_0.pc_nxt_14_ )
  );
  NOR2X1 _10970_ (
    .A(_03795_),
    .B( execution_unit_0.pc_sw_15_ ),
    .Y(_03651_)
  );
  OAI21X1 _10971_ (
    .A(_03811_),
    .B(_03643_),
    .C(_03812_),
    .Y(_03652_)
  );
  NAND3X1 _10972_ (
    .A( dbg_0.UNUSED_pc_14_ ),
    .B( dbg_0.UNUSED_pc_15_ ),
    .C(_03642_),
    .Y(_03653_)
  );
  NAND3X1 _10973_ (
    .A(_03547_),
    .B(_03652_),
    .C(_03653_),
    .Y(_03654_)
  );
  AOI21X1 _10974_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03546_),
    .C(_03564_),
    .Y(_03655_)
  );
  AOI21X1 _10975_ (
    .A(_03654_),
    .B(_03655_),
    .C(_03651_),
    .Y( execution_unit_0.pc_nxt_15_ )
  );
  NOR2X1 _10976_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03656_)
  );
  NAND2X1 _10977_ (
    .A(_03761_),
    .B(_03656_),
    .Y(_03657_)
  );
  OR2X1 _10978_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03657_),
    .Y(_03658_)
  );
  NOR2X1 _10979_ (
    .A( execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03555_),
    .Y(_03659_)
  );
  OR2X1 _10980_ (
    .A( execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03555_),
    .Y(_03660_)
  );
  NOR2X1 _10981_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( dbg_0.cpu_stat_full_0_ ),
    .Y(_03661_)
  );
  OAI21X1 _10982_ (
    .A(_03658_),
    .B(_03660_),
    .C(_03661_),
    .Y(_03662_)
  );
  NAND2X1 _10983_ (
    .A(_03814_),
    .B(_03815_),
    .Y(_03663_)
  );
  OR2X1 _10984_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_03663_),
    .Y(_03664_)
  );
  OAI21X1 _10985_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_03664_),
    .C( dbg_0.cpu_stat_full_0_ ),
    .Y(_03665_)
  );
  AND2X1 _10986_ (
    .A(_03662_),
    .B(_03665_),
    .Y( execution_unit_0.inst_dest_0_ )
  );
  AND2X1 _10987_ (
    .A(_03763_),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03666_)
  );
  NAND2X1 _10988_ (
    .A(_03761_),
    .B(_03666_),
    .Y(_03667_)
  );
  NOR2X1 _10989_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03667_),
    .Y(_03668_)
  );
  OAI21X1 _10990_ (
    .A(_03660_),
    .B(_03668_),
    .C(_03661_),
    .Y(_03669_)
  );
  NAND3X1 _10991_ (
    .A(_03813_),
    .B(_03814_),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03670_)
  );
  XOR2X1 _10992_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_03664_),
    .Y(_03671_)
  );
  NAND2X1 _10993_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_03671_),
    .Y(_03672_)
  );
  OAI21X1 _10994_ (
    .A(_03670_),
    .B(_03672_),
    .C(_03669_),
    .Y( execution_unit_0.inst_dest_1_ )
  );
  NOR2X1 _10995_ (
    .A(_03763_),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03673_)
  );
  NAND2X1 _10996_ (
    .A(_03761_),
    .B(_03673_),
    .Y(_03674_)
  );
  OR2X1 _10997_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03674_),
    .Y(_03675_)
  );
  NAND2X1 _10998_ (
    .A(_03659_),
    .B(_03661_),
    .Y(_03676_)
  );
  NAND3X1 _10999_ (
    .A(_03813_),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C(_03815_),
    .Y(_03677_)
  );
  OAI22X1 _11000_ (
    .A(_03675_),
    .B(_03676_),
    .C(_03677_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_2_ )
  );
  NAND2X1 _11001_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03678_)
  );
  NOR2X1 _11002_ (
    .A( frontend_0.inst_dest_bin_2_ ),
    .B(_03678_),
    .Y(_03679_)
  );
  NAND2X1 _11003_ (
    .A(_03760_),
    .B(_03679_),
    .Y(_03680_)
  );
  NAND3X1 _11004_ (
    .A(_03813_),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03681_)
  );
  OAI22X1 _11005_ (
    .A(_03676_),
    .B(_03680_),
    .C(_03681_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_3_ )
  );
  NAND3X1 _11006_ (
    .A(_03760_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03656_),
    .Y(_03682_)
  );
  OR2X1 _11007_ (
    .A(_03813_),
    .B(_03663_),
    .Y(_03683_)
  );
  OAI22X1 _11008_ (
    .A(_03676_),
    .B(_03682_),
    .C(_03683_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_4_ )
  );
  NAND3X1 _11009_ (
    .A(_03760_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03666_),
    .Y(_03684_)
  );
  NAND3X1 _11010_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_03814_),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03685_)
  );
  OAI22X1 _11011_ (
    .A(_03676_),
    .B(_03684_),
    .C(_03685_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_5_ )
  );
  NAND3X1 _11012_ (
    .A(_03760_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03673_),
    .Y(_03686_)
  );
  NAND3X1 _11013_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C(_03815_),
    .Y(_03687_)
  );
  OAI22X1 _11014_ (
    .A(_03676_),
    .B(_03686_),
    .C(_03687_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_6_ )
  );
  OR2X1 _11015_ (
    .A(_03761_),
    .B(_03678_),
    .Y(_03688_)
  );
  OR2X1 _11016_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03688_),
    .Y(_03689_)
  );
  NAND3X1 _11017_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03690_)
  );
  OAI22X1 _11018_ (
    .A(_03676_),
    .B(_03689_),
    .C(_03690_),
    .D(_03672_),
    .Y( execution_unit_0.inst_dest_7_ )
  );
  OR2X1 _11019_ (
    .A(_03760_),
    .B(_03657_),
    .Y(_03691_)
  );
  OAI22X1 _11020_ (
    .A(_03664_),
    .B(_03665_),
    .C(_03676_),
    .D(_03691_),
    .Y( execution_unit_0.inst_dest_8_ )
  );
  OR2X1 _11021_ (
    .A(_03760_),
    .B(_03667_),
    .Y(_03692_)
  );
  OR2X1 _11022_ (
    .A(_03786_),
    .B(_03671_),
    .Y(_03693_)
  );
  OAI22X1 _11023_ (
    .A(_03676_),
    .B(_03692_),
    .C(_03693_),
    .D(_03670_),
    .Y( execution_unit_0.inst_dest_9_ )
  );
  OR2X1 _11024_ (
    .A(_03760_),
    .B(_03674_),
    .Y(_03694_)
  );
  OAI22X1 _11025_ (
    .A(_03677_),
    .B(_03693_),
    .C(_03694_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_10_ )
  );
  NAND2X1 _11026_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03679_),
    .Y(_03695_)
  );
  OAI22X1 _11027_ (
    .A(_03681_),
    .B(_03693_),
    .C(_03695_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_11_ )
  );
  NAND3X1 _11028_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03656_),
    .Y(_03696_)
  );
  OAI22X1 _11029_ (
    .A(_03683_),
    .B(_03693_),
    .C(_03696_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_12_ )
  );
  NAND3X1 _11030_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03666_),
    .Y(_03697_)
  );
  OAI22X1 _11031_ (
    .A(_03685_),
    .B(_03693_),
    .C(_03697_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_13_ )
  );
  NAND3X1 _11032_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03673_),
    .Y(_03698_)
  );
  OAI22X1 _11033_ (
    .A(_03687_),
    .B(_03693_),
    .C(_03698_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_14_ )
  );
  OR2X1 _11034_ (
    .A(_03760_),
    .B(_03688_),
    .Y(_03699_)
  );
  OAI22X1 _11035_ (
    .A(_03690_),
    .B(_03693_),
    .C(_03699_),
    .D(_03676_),
    .Y( execution_unit_0.inst_dest_15_ )
  );
  OAI21X1 _11036_ (
    .A(_03754_),
    .B(_03658_),
    .C(_03755_),
    .Y(_03700_)
  );
  NOR2X1 _11037_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_03701_)
  );
  NAND2X1 _11038_ (
    .A(_03700_),
    .B(_03701_),
    .Y(_03702_)
  );
  NAND2X1 _11039_ (
    .A(_03765_),
    .B(_03767_),
    .Y(_03703_)
  );
  OR2X1 _11040_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03703_),
    .Y(_03704_)
  );
  OR2X1 _11041_ (
    .A( frontend_0.inst_jmp_bin_1_ ),
    .B(_03704_),
    .Y(_03705_)
  );
  OAI21X1 _11042_ (
    .A(_03752_),
    .B(_03705_),
    .C(_03702_),
    .Y( execution_unit_0.inst_src_0_ )
  );
  NOR2X1 _11043_ (
    .A(_03754_),
    .B( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_03706_)
  );
  AOI21X1 _11044_ (
    .A(_03668_),
    .B(_03706_),
    .C( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_03707_)
  );
  NAND3X1 _11045_ (
    .A(_03758_),
    .B(_03765_),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03708_)
  );
  XOR2X1 _11046_ (
    .A( frontend_0.inst_jmp_bin_1_ ),
    .B(_03704_),
    .Y(_03709_)
  );
  NAND2X1 _11047_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B(_03709_),
    .Y(_03710_)
  );
  OAI22X1 _11048_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B(_03707_),
    .C(_03708_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_1_ )
  );
  NAND2X1 _11049_ (
    .A(_03701_),
    .B(_03706_),
    .Y(_03711_)
  );
  NAND3X1 _11050_ (
    .A(_03758_),
    .B( frontend_0.inst_src_bin_1_ ),
    .C(_03767_),
    .Y(_03712_)
  );
  OAI22X1 _11051_ (
    .A(_03675_),
    .B(_03711_),
    .C(_03712_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_2_ )
  );
  NAND3X1 _11052_ (
    .A(_03758_),
    .B( frontend_0.inst_src_bin_1_ ),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03713_)
  );
  OAI22X1 _11053_ (
    .A(_03680_),
    .B(_03711_),
    .C(_03713_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_3_ )
  );
  OR2X1 _11054_ (
    .A(_03758_),
    .B(_03703_),
    .Y(_03714_)
  );
  OAI22X1 _11055_ (
    .A(_03682_),
    .B(_03711_),
    .C(_03714_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_4_ )
  );
  NAND3X1 _11056_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03765_),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03715_)
  );
  OAI22X1 _11057_ (
    .A(_03684_),
    .B(_03711_),
    .C(_03715_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_5_ )
  );
  NAND3X1 _11058_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B( frontend_0.inst_src_bin_1_ ),
    .C(_03767_),
    .Y(_03716_)
  );
  OAI22X1 _11059_ (
    .A(_03686_),
    .B(_03711_),
    .C(_03716_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_6_ )
  );
  NAND3X1 _11060_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B( frontend_0.inst_src_bin_1_ ),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03717_)
  );
  OAI22X1 _11061_ (
    .A(_03689_),
    .B(_03711_),
    .C(_03717_),
    .D(_03710_),
    .Y( execution_unit_0.inst_src_7_ )
  );
  NAND2X1 _11062_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .Y(_03718_)
  );
  OAI22X1 _11063_ (
    .A(_03691_),
    .B(_03711_),
    .C(_03718_),
    .D(_03704_),
    .Y( execution_unit_0.inst_src_8_ )
  );
  OR2X1 _11064_ (
    .A(_03752_),
    .B(_03709_),
    .Y(_03719_)
  );
  OAI22X1 _11065_ (
    .A(_03692_),
    .B(_03711_),
    .C(_03719_),
    .D(_03708_),
    .Y( execution_unit_0.inst_src_9_ )
  );
  OAI22X1 _11066_ (
    .A(_03694_),
    .B(_03711_),
    .C(_03712_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_10_ )
  );
  OAI22X1 _11067_ (
    .A(_03695_),
    .B(_03711_),
    .C(_03713_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_11_ )
  );
  OAI22X1 _11068_ (
    .A(_03696_),
    .B(_03711_),
    .C(_03714_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_12_ )
  );
  OAI22X1 _11069_ (
    .A(_03697_),
    .B(_03711_),
    .C(_03715_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_13_ )
  );
  OAI22X1 _11070_ (
    .A(_03698_),
    .B(_03711_),
    .C(_03716_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_14_ )
  );
  OAI22X1 _11071_ (
    .A(_03699_),
    .B(_03711_),
    .C(_03717_),
    .D(_03719_),
    .Y( execution_unit_0.inst_src_15_ )
  );
  NAND2X1 _11072_ (
    .A(_03744_),
    .B(_03745_),
    .Y(_03720_)
  );
  OR2X1 _11073_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03720_),
    .Y(_03721_)
  );
  OR2X1 _11074_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03721_),
    .Y(_03722_)
  );
  NOR2X1 _11075_ (
    .A(_03538_),
    .B(_03722_),
    .Y(_06248_)
  );
  NAND3X1 _11076_ (
    .A(_03743_),
    .B(_03744_),
    .C( frontend_0.irq_addr_1_ ),
    .Y(_03723_)
  );
  XOR2X1 _11077_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03721_),
    .Y(_03724_)
  );
  NAND2X1 _11078_ (
    .A(_03537_),
    .B(_03724_),
    .Y(_03725_)
  );
  NOR2X1 _11079_ (
    .A(_03723_),
    .B(_03725_),
    .Y(_06253_)
  );
  NAND3X1 _11080_ (
    .A(_03743_),
    .B( frontend_0.irq_addr_2_ ),
    .C(_03745_),
    .Y(_03726_)
  );
  NOR2X1 _11081_ (
    .A(_03725_),
    .B(_03726_),
    .Y(_06254_)
  );
  NAND2X1 _11082_ (
    .A( frontend_0.irq_addr_2_ ),
    .B( frontend_0.irq_addr_1_ ),
    .Y(_03727_)
  );
  OR2X1 _11083_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03727_),
    .Y(_03728_)
  );
  NOR2X1 _11084_ (
    .A(_03725_),
    .B(_03728_),
    .Y(_06255_)
  );
  OR2X1 _11085_ (
    .A(_03743_),
    .B(_03720_),
    .Y(_03729_)
  );
  NOR2X1 _11086_ (
    .A(_03725_),
    .B(_03729_),
    .Y(_06256_)
  );
  NAND3X1 _11087_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03744_),
    .C( frontend_0.irq_addr_1_ ),
    .Y(_03730_)
  );
  NOR2X1 _11088_ (
    .A(_03725_),
    .B(_03730_),
    .Y(_06257_)
  );
  NAND3X1 _11089_ (
    .A( frontend_0.irq_addr_3_ ),
    .B( frontend_0.irq_addr_2_ ),
    .C(_03745_),
    .Y(_03731_)
  );
  NOR2X1 _11090_ (
    .A(_03725_),
    .B(_03731_),
    .Y(_06258_)
  );
  NAND3X1 _11091_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03537_),
    .C(_03724_),
    .Y(_03732_)
  );
  NOR2X1 _11092_ (
    .A(_03727_),
    .B(_03732_),
    .Y(_06259_)
  );
  NOR2X1 _11093_ (
    .A(_03596_),
    .B(_03721_),
    .Y(_06260_)
  );
  OR2X1 _11094_ (
    .A(_03538_),
    .B(_03724_),
    .Y(_03733_)
  );
  NOR2X1 _11095_ (
    .A(_03723_),
    .B(_03733_),
    .Y(_06261_)
  );
  NOR2X1 _11096_ (
    .A(_03726_),
    .B(_03733_),
    .Y(_06249_)
  );
  NOR2X1 _11097_ (
    .A(_03728_),
    .B(_03733_),
    .Y(_06250_)
  );
  NOR2X1 _11098_ (
    .A(_03596_),
    .B(_03729_),
    .Y(_06251_)
  );
  NOR2X1 _11099_ (
    .A(_03730_),
    .B(_03733_),
    .Y(_06252_)
  );
  OAI21X1 _11100_ (
    .A(_03786_),
    .B(_03855_),
    .C(_03816_),
    .Y(_03734_)
  );
  NOR2X1 _11101_ (
    .A(_03564_),
    .B(_03734_),
    .Y(_03735_)
  );
  OAI21X1 _11102_ (
    .A(_03568_),
    .B(_03570_),
    .C(_03735_),
    .Y( frontend_0.mb_en )
  );
  NAND2X1 _11103_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_03758_),
    .Y(_03736_)
  );
  OR2X1 _11104_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .Y(_03737_)
  );
  NOR2X1 _11105_ (
    .A(_03736_),
    .B(_03737_),
    .Y( execution_unit_0.alu_0.inst_jmp_0_ )
  );
  NAND2X1 _11106_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( frontend_0.inst_jmp_bin_0_ ),
    .Y(_03738_)
  );
  NOR2X1 _11107_ (
    .A(_03737_),
    .B(_03738_),
    .Y( execution_unit_0.alu_0.inst_jmp_1_ )
  );
  NAND3X1 _11108_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .C(_03758_),
    .Y(_03739_)
  );
  NOR2X1 _11109_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03739_),
    .Y( execution_unit_0.alu_0.inst_jmp_2_ )
  );
  NAND3X1 _11110_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .C( frontend_0.inst_jmp_bin_0_ ),
    .Y(_03740_)
  );
  NOR2X1 _11111_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03740_),
    .Y( execution_unit_0.alu_0.inst_jmp_3_ )
  );
  OR2X1 _11112_ (
    .A(_03757_),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .Y(_03741_)
  );
  NOR2X1 _11113_ (
    .A(_03736_),
    .B(_03741_),
    .Y( execution_unit_0.alu_0.inst_jmp_4_ )
  );
  NOR2X1 _11114_ (
    .A(_03738_),
    .B(_03741_),
    .Y( execution_unit_0.alu_0.inst_jmp_5_ )
  );
  NOR2X1 _11115_ (
    .A(_03757_),
    .B(_03739_),
    .Y( execution_unit_0.alu_0.inst_jmp_6_ )
  );
  NAND3X1 _11116_ (
    .A(_03855_),
    .B( frontend_0.i_state_nxt_0_ ),
    .C( frontend_0.i_state_nxt_2_ ),
    .Y(_03742_)
  );
  INVX1 _11117_ (
    .A(_03742_),
    .Y(_03253_)
  );
  INVX1 _11118_ (
    .A(_06327_),
    .Y(_03255_)
  );
  INVX1 _11119_ (
    .A(_06327_),
    .Y(_03256_)
  );
  INVX1 _11120_ (
    .A(_06327_),
    .Y(_03257_)
  );
  INVX1 _11121_ (
    .A(_06327_),
    .Y(_03258_)
  );
  INVX1 _11122_ (
    .A(_06327_),
    .Y(_03259_)
  );
  INVX1 _11123_ (
    .A(_06327_),
    .Y(_03260_)
  );
  INVX1 _11124_ (
    .A(_06327_),
    .Y(_03261_)
  );
  INVX1 _11125_ (
    .A(_06327_),
    .Y(_03262_)
  );
  INVX1 _11126_ (
    .A(_06327_),
    .Y(_03263_)
  );
  INVX1 _11127_ (
    .A(_06327_),
    .Y(_03264_)
  );
  INVX1 _11128_ (
    .A(_06327_),
    .Y(_03265_)
  );
  INVX1 _11129_ (
    .A(_06327_),
    .Y(_03266_)
  );
  INVX1 _11130_ (
    .A(_06327_),
    .Y(_03267_)
  );
  INVX1 _11131_ (
    .A(_06327_),
    .Y(_03268_)
  );
  INVX1 _11132_ (
    .A(_06327_),
    .Y(_03269_)
  );
  INVX1 _11133_ (
    .A(_06327_),
    .Y(_03270_)
  );
  INVX1 _11134_ (
    .A(_06327_),
    .Y(_03271_)
  );
  INVX1 _11135_ (
    .A(_06327_),
    .Y(_03272_)
  );
  INVX1 _11136_ (
    .A(_06327_),
    .Y(_03273_)
  );
  INVX1 _11137_ (
    .A(_06327_),
    .Y(_03274_)
  );
  INVX1 _11138_ (
    .A(_06327_),
    .Y(_03275_)
  );
  INVX1 _11139_ (
    .A(_06327_),
    .Y(_03276_)
  );
  INVX1 _11140_ (
    .A(_06327_),
    .Y(_03277_)
  );
  INVX1 _11141_ (
    .A(_06327_),
    .Y(_03278_)
  );
  INVX1 _11142_ (
    .A(_06327_),
    .Y(_03279_)
  );
  INVX1 _11143_ (
    .A(_06327_),
    .Y(_03280_)
  );
  INVX1 _11144_ (
    .A(_06327_),
    .Y(_03281_)
  );
  INVX1 _11145_ (
    .A(_06327_),
    .Y(_03282_)
  );
  INVX1 _11146_ (
    .A(_06327_),
    .Y(_03283_)
  );
  INVX1 _11147_ (
    .A(_06327_),
    .Y(_03284_)
  );
  INVX1 _11148_ (
    .A(_06327_),
    .Y(_03285_)
  );
  INVX1 _11149_ (
    .A(_06327_),
    .Y(_03286_)
  );
  INVX1 _11150_ (
    .A(_06327_),
    .Y(_03287_)
  );
  INVX1 _11151_ (
    .A(_06327_),
    .Y(_03288_)
  );
  INVX1 _11152_ (
    .A(_06327_),
    .Y(_03289_)
  );
  INVX1 _11153_ (
    .A(_06327_),
    .Y(_03290_)
  );
  INVX1 _11154_ (
    .A(_06327_),
    .Y(_03291_)
  );
  INVX1 _11155_ (
    .A(_06327_),
    .Y(_03292_)
  );
  INVX1 _11156_ (
    .A(_06327_),
    .Y(_03293_)
  );
  INVX1 _11157_ (
    .A(_06327_),
    .Y(_03294_)
  );
  INVX1 _11158_ (
    .A(_06327_),
    .Y(_03295_)
  );
  INVX1 _11159_ (
    .A(_06327_),
    .Y(_03296_)
  );
  INVX1 _11160_ (
    .A(_06327_),
    .Y(_03297_)
  );
  INVX1 _11161_ (
    .A(_06327_),
    .Y(_03298_)
  );
  INVX1 _11162_ (
    .A(_06327_),
    .Y(_03299_)
  );
  INVX1 _11163_ (
    .A(_06327_),
    .Y(_03300_)
  );
  INVX1 _11164_ (
    .A(_06327_),
    .Y(_03301_)
  );
  INVX1 _11165_ (
    .A(_06327_),
    .Y(_03302_)
  );
  INVX1 _11166_ (
    .A(_06327_),
    .Y(_03303_)
  );
  INVX1 _11167_ (
    .A(_06327_),
    .Y(_03304_)
  );
  INVX1 _11168_ (
    .A(_06327_),
    .Y(_03305_)
  );
  INVX1 _11169_ (
    .A(_06327_),
    .Y(_03306_)
  );
  INVX1 _11170_ (
    .A(_06327_),
    .Y(_03307_)
  );
  INVX1 _11171_ (
    .A(_06327_),
    .Y(_03308_)
  );
  INVX1 _11172_ (
    .A(_06327_),
    .Y(_03309_)
  );
  INVX1 _11173_ (
    .A(_06327_),
    .Y(_03310_)
  );
  INVX1 _11174_ (
    .A(_06327_),
    .Y(_03311_)
  );
  INVX1 _11175_ (
    .A(_06327_),
    .Y(_03312_)
  );
  INVX1 _11176_ (
    .A(_06327_),
    .Y(_03313_)
  );
  INVX1 _11177_ (
    .A(_06327_),
    .Y(_03314_)
  );
  INVX1 _11178_ (
    .A(_06327_),
    .Y(_03315_)
  );
  INVX1 _11179_ (
    .A(_06327_),
    .Y(_03316_)
  );
  INVX1 _11180_ (
    .A(_06327_),
    .Y(_03317_)
  );
  INVX1 _11181_ (
    .A(_06327_),
    .Y(_03318_)
  );
  INVX1 _11182_ (
    .A(_06327_),
    .Y(_03319_)
  );
  INVX1 _11183_ (
    .A(_06327_),
    .Y(_03320_)
  );
  INVX1 _11184_ (
    .A(_06327_),
    .Y(_03321_)
  );
  INVX1 _11185_ (
    .A(_06327_),
    .Y(_03322_)
  );
  INVX1 _11186_ (
    .A(_06327_),
    .Y(_03323_)
  );
  INVX1 _11187_ (
    .A(_06327_),
    .Y(_03324_)
  );
  INVX1 _11188_ (
    .A(_06327_),
    .Y(_03325_)
  );
  INVX1 _11189_ (
    .A(_06327_),
    .Y(_03326_)
  );
  INVX1 _11190_ (
    .A(_06327_),
    .Y(_03327_)
  );
  INVX1 _11191_ (
    .A(_06327_),
    .Y(_03328_)
  );
  INVX1 _11192_ (
    .A(_06327_),
    .Y(_03329_)
  );
  INVX1 _11193_ (
    .A(_06327_),
    .Y(_03330_)
  );
  INVX1 _11194_ (
    .A(_06327_),
    .Y(_03331_)
  );
  INVX1 _11195_ (
    .A(_06327_),
    .Y(_03332_)
  );
  INVX1 _11196_ (
    .A(_06327_),
    .Y(_03333_)
  );
  INVX1 _11197_ (
    .A(_06327_),
    .Y(_03334_)
  );
  INVX1 _11198_ (
    .A(_06327_),
    .Y(_03335_)
  );
  INVX1 _11199_ (
    .A(_06327_),
    .Y(_03336_)
  );
  INVX1 _11200_ (
    .A(_06327_),
    .Y(_03337_)
  );
  INVX1 _11201_ (
    .A(_06327_),
    .Y(_03338_)
  );
  INVX1 _11202_ (
    .A(_06327_),
    .Y(_03339_)
  );
  INVX1 _11203_ (
    .A(_06327_),
    .Y(_03340_)
  );
  INVX1 _11204_ (
    .A(_06327_),
    .Y(_03341_)
  );
  INVX1 _11205_ (
    .A(_06327_),
    .Y(_03342_)
  );
  INVX1 _11206_ (
    .A(_06327_),
    .Y(_03343_)
  );
  INVX1 _11207_ (
    .A(_06327_),
    .Y(_03344_)
  );
  INVX1 _11208_ (
    .A(_06327_),
    .Y(_03345_)
  );
  INVX1 _11209_ (
    .A(_06327_),
    .Y(_03346_)
  );
  INVX1 _11210_ (
    .A(_06327_),
    .Y(_03347_)
  );
  INVX1 _11211_ (
    .A(_06327_),
    .Y(_03348_)
  );
  INVX1 _11212_ (
    .A(_06327_),
    .Y(_03349_)
  );
  INVX1 _11213_ (
    .A(_06327_),
    .Y(_03350_)
  );
  INVX1 _11214_ (
    .A(_06327_),
    .Y(_03351_)
  );
  INVX1 _11215_ (
    .A(_06327_),
    .Y(_03352_)
  );
  INVX1 _11216_ (
    .A(_06327_),
    .Y(_03353_)
  );
  INVX1 _11217_ (
    .A(_06327_),
    .Y(_03354_)
  );
  INVX1 _11218_ (
    .A(_06327_),
    .Y(_03355_)
  );
  INVX1 _11219_ (
    .A(_06327_),
    .Y(_03356_)
  );
  INVX1 _11220_ (
    .A(_06327_),
    .Y(_03357_)
  );
  INVX1 _11221_ (
    .A(_06327_),
    .Y(_03358_)
  );
  INVX1 _11222_ (
    .A(_06327_),
    .Y(_03359_)
  );
  INVX1 _11223_ (
    .A(_06327_),
    .Y(_03360_)
  );
  INVX1 _11224_ (
    .A(_06327_),
    .Y(_03361_)
  );
  INVX1 _11225_ (
    .A(_06327_),
    .Y(_03362_)
  );
  INVX1 _11226_ (
    .A(_06327_),
    .Y(_03363_)
  );
  INVX1 _11227_ (
    .A(_06327_),
    .Y(_03364_)
  );
  INVX1 _11228_ (
    .A(_06327_),
    .Y(_03365_)
  );
  INVX1 _11229_ (
    .A(_06327_),
    .Y(_03366_)
  );
  DFFSR _11230_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_0_ ),
    .Q( execution_unit_0.e_state_0_ ),
    .R(1'h1),
    .S(_03254_)
  );
  DFFSR _11231_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_1_ ),
    .Q( execution_unit_0.e_state_1_ ),
    .R(_03255_),
    .S(1'h1)
  );
  DFFSR _11232_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_2_ ),
    .Q( execution_unit_0.e_state_2_ ),
    .R(_03256_),
    .S(1'h1)
  );
  DFFSR _11233_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_3_ ),
    .Q( execution_unit_0.e_state_3_ ),
    .R(_03257_),
    .S(1'h1)
  );
  DFFSR _11234_ (
    .CLK(dco_clk),
    .D(_03367_),
    .Q( execution_unit_0.alu_0.inst_alu_0_ ),
    .R(_03258_),
    .S(1'h1)
  );
  DFFSR _11235_ (
    .CLK(dco_clk),
    .D(_03368_),
    .Q( execution_unit_0.alu_0.inst_alu_1_ ),
    .R(_03259_),
    .S(1'h1)
  );
  DFFSR _11236_ (
    .CLK(dco_clk),
    .D(_03369_),
    .Q( execution_unit_0.alu_0.inst_alu_2_ ),
    .R(_03260_),
    .S(1'h1)
  );
  DFFSR _11237_ (
    .CLK(dco_clk),
    .D(_03370_),
    .Q( execution_unit_0.alu_0.inst_alu_3_ ),
    .R(_03261_),
    .S(1'h1)
  );
  DFFSR _11238_ (
    .CLK(dco_clk),
    .D(_03371_),
    .Q( execution_unit_0.alu_0.inst_alu_4_ ),
    .R(_03262_),
    .S(1'h1)
  );
  DFFSR _11239_ (
    .CLK(dco_clk),
    .D(_03372_),
    .Q( execution_unit_0.alu_0.inst_alu_5_ ),
    .R(_03263_),
    .S(1'h1)
  );
  DFFSR _11240_ (
    .CLK(dco_clk),
    .D(_03373_),
    .Q( execution_unit_0.alu_0.inst_alu_6_ ),
    .R(_03264_),
    .S(1'h1)
  );
  DFFSR _11241_ (
    .CLK(dco_clk),
    .D(_03374_),
    .Q( execution_unit_0.alu_0.inst_alu_7_ ),
    .R(_03265_),
    .S(1'h1)
  );
  DFFSR _11242_ (
    .CLK(dco_clk),
    .D(_03375_),
    .Q( execution_unit_0.alu_0.inst_alu_8_ ),
    .R(_03266_),
    .S(1'h1)
  );
  DFFSR _11243_ (
    .CLK(dco_clk),
    .D(_03376_),
    .Q( execution_unit_0.alu_0.inst_alu_9_ ),
    .R(_03267_),
    .S(1'h1)
  );
  DFFSR _11244_ (
    .CLK(dco_clk),
    .D(_03377_),
    .Q( execution_unit_0.alu_0.inst_alu_10_ ),
    .R(_03268_),
    .S(1'h1)
  );
  DFFSR _11245_ (
    .CLK(dco_clk),
    .D(_03378_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .R(_03269_),
    .S(1'h1)
  );
  DFFSR _11246_ (
    .CLK(dco_clk),
    .D(_03379_),
    .Q( frontend_0.exec_dext_rdy ),
    .R(_03270_),
    .S(1'h1)
  );
  DFFSR _11247_ (
    .CLK(dco_clk),
    .D(_03380_),
    .Q( frontend_0.exec_src_wr ),
    .R(_03271_),
    .S(1'h1)
  );
  DFFSR _11248_ (
    .CLK(dco_clk),
    .D(_03381_),
    .Q( frontend_0.exec_dst_wr ),
    .R(_03272_),
    .S(1'h1)
  );
  DFFSR _11249_ (
    .CLK(dco_clk),
    .D(_03382_),
    .Q( frontend_0.exec_jmp ),
    .R(_03273_),
    .S(1'h1)
  );
  DFFSR _11250_ (
    .CLK(dco_clk),
    .D(_03383_),
    .Q( frontend_0.inst_sz_0_ ),
    .R(_03274_),
    .S(1'h1)
  );
  DFFSR _11251_ (
    .CLK(dco_clk),
    .D(_03384_),
    .Q( frontend_0.inst_sz_1_ ),
    .R(_03275_),
    .S(1'h1)
  );
  DFFSR _11252_ (
    .CLK(dco_clk),
    .D(_03385_),
    .Q( execution_unit_0.alu_0.inst_bw ),
    .R(_03276_),
    .S(1'h1)
  );
  DFFSR _11253_ (
    .CLK(dco_clk),
    .D(_03386_),
    .Q( execution_unit_0.inst_as_0_ ),
    .R(_03277_),
    .S(1'h1)
  );
  DFFSR _11254_ (
    .CLK(dco_clk),
    .D(_03387_),
    .Q( execution_unit_0.inst_as_1_ ),
    .R(_03278_),
    .S(1'h1)
  );
  DFFSR _11255_ (
    .CLK(dco_clk),
    .D(_03388_),
    .Q( execution_unit_0.inst_as_2_ ),
    .R(_03279_),
    .S(1'h1)
  );
  DFFSR _11256_ (
    .CLK(dco_clk),
    .D(_03389_),
    .Q( execution_unit_0.inst_as_3_ ),
    .R(_03280_),
    .S(1'h1)
  );
  DFFSR _11257_ (
    .CLK(dco_clk),
    .D(_03390_),
    .Q( execution_unit_0.inst_as_4_ ),
    .R(_03281_),
    .S(1'h1)
  );
  DFFSR _11258_ (
    .CLK(dco_clk),
    .D(_03391_),
    .Q( execution_unit_0.inst_as_5_ ),
    .R(_03282_),
    .S(1'h1)
  );
  DFFSR _11259_ (
    .CLK(dco_clk),
    .D(_03392_),
    .Q( execution_unit_0.inst_as_6_ ),
    .R(_03283_),
    .S(1'h1)
  );
  DFFSR _11260_ (
    .CLK(dco_clk),
    .D(_03393_),
    .Q( execution_unit_0.inst_as_7_ ),
    .R(_03284_),
    .S(1'h1)
  );
  DFFSR _11261_ (
    .CLK(dco_clk),
    .D(_03394_),
    .Q( frontend_0.inst_src_bin_0_ ),
    .R(_03285_),
    .S(1'h1)
  );
  DFFSR _11262_ (
    .CLK(dco_clk),
    .D(_03395_),
    .Q( frontend_0.inst_src_bin_1_ ),
    .R(_03286_),
    .S(1'h1)
  );
  DFFSR _11263_ (
    .CLK(dco_clk),
    .D(_03396_),
    .Q( frontend_0.inst_dest_bin_0_ ),
    .R(_03287_),
    .S(1'h1)
  );
  DFFSR _11264_ (
    .CLK(dco_clk),
    .D(_03397_),
    .Q( frontend_0.inst_dest_bin_1_ ),
    .R(_03288_),
    .S(1'h1)
  );
  DFFSR _11265_ (
    .CLK(dco_clk),
    .D(_03398_),
    .Q( frontend_0.inst_dest_bin_2_ ),
    .R(_03289_),
    .S(1'h1)
  );
  DFFSR _11266_ (
    .CLK(dco_clk),
    .D(_03399_),
    .Q( frontend_0.inst_dest_bin_3_ ),
    .R(_03290_),
    .S(1'h1)
  );
  DFFSR _11267_ (
    .CLK(dco_clk),
    .D(_03400_),
    .Q( execution_unit_0.inst_mov ),
    .R(_03291_),
    .S(1'h1)
  );
  DFFSR _11268_ (
    .CLK(dco_clk),
    .D(_03401_),
    .Q( frontend_0.inst_jmp_bin_0_ ),
    .R(_03292_),
    .S(1'h1)
  );
  DFFSR _11269_ (
    .CLK(dco_clk),
    .D(_03402_),
    .Q( frontend_0.inst_jmp_bin_1_ ),
    .R(_03293_),
    .S(1'h1)
  );
  DFFSR _11270_ (
    .CLK(dco_clk),
    .D(_03403_),
    .Q( frontend_0.inst_jmp_bin_2_ ),
    .R(_03294_),
    .S(1'h1)
  );
  DFFSR _11271_ (
    .CLK(dco_clk),
    .D(_03404_),
    .Q( execution_unit_0.alu_0.inst_so_0_ ),
    .R(_03295_),
    .S(1'h1)
  );
  DFFSR _11272_ (
    .CLK(dco_clk),
    .D(_03405_),
    .Q( execution_unit_0.alu_0.inst_so_1_ ),
    .R(_03296_),
    .S(1'h1)
  );
  DFFSR _11273_ (
    .CLK(dco_clk),
    .D(_03406_),
    .Q( execution_unit_0.alu_0.inst_so_3_ ),
    .R(_03297_),
    .S(1'h1)
  );
  DFFSR _11274_ (
    .CLK(dco_clk),
    .D(_03407_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .R(_03298_),
    .S(1'h1)
  );
  DFFSR _11275_ (
    .CLK(dco_clk),
    .D(_03408_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .R(_03299_),
    .S(1'h1)
  );
  DFFSR _11276_ (
    .CLK(dco_clk),
    .D(_03409_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .R(_03300_),
    .S(1'h1)
  );
  DFFSR _11277_ (
    .CLK(dco_clk),
    .D(_03410_),
    .Q( execution_unit_0.alu_0.inst_so_7_ ),
    .R(_03301_),
    .S(1'h1)
  );
  DFFSR _11278_ (
    .CLK(dco_clk),
    .D(_03411_),
    .Q( execution_unit_0.inst_type_0_ ),
    .R(_03302_),
    .S(1'h1)
  );
  DFFSR _11279_ (
    .CLK(dco_clk),
    .D(_03412_),
    .Q( execution_unit_0.inst_type_1_ ),
    .R(_03303_),
    .S(1'h1)
  );
  DFFSR _11280_ (
    .CLK(dco_clk),
    .D(_03413_),
    .Q( execution_unit_0.inst_type_2_ ),
    .R(_03304_),
    .S(1'h1)
  );
  DFFSR _11281_ (
    .CLK(dco_clk),
    .D(_03414_),
    .Q( execution_unit_0.inst_dext_0_ ),
    .R(_03305_),
    .S(1'h1)
  );
  DFFSR _11282_ (
    .CLK(dco_clk),
    .D(_03415_),
    .Q( execution_unit_0.inst_dext_1_ ),
    .R(_03306_),
    .S(1'h1)
  );
  DFFSR _11283_ (
    .CLK(dco_clk),
    .D(_03416_),
    .Q( execution_unit_0.inst_dext_2_ ),
    .R(_03307_),
    .S(1'h1)
  );
  DFFSR _11284_ (
    .CLK(dco_clk),
    .D(_03417_),
    .Q( execution_unit_0.inst_dext_3_ ),
    .R(_03308_),
    .S(1'h1)
  );
  DFFSR _11285_ (
    .CLK(dco_clk),
    .D(_03418_),
    .Q( execution_unit_0.inst_dext_4_ ),
    .R(_03309_),
    .S(1'h1)
  );
  DFFSR _11286_ (
    .CLK(dco_clk),
    .D(_03419_),
    .Q( execution_unit_0.inst_dext_5_ ),
    .R(_03310_),
    .S(1'h1)
  );
  DFFSR _11287_ (
    .CLK(dco_clk),
    .D(_03420_),
    .Q( execution_unit_0.inst_dext_6_ ),
    .R(_03311_),
    .S(1'h1)
  );
  DFFSR _11288_ (
    .CLK(dco_clk),
    .D(_03421_),
    .Q( execution_unit_0.inst_dext_7_ ),
    .R(_03312_),
    .S(1'h1)
  );
  DFFSR _11289_ (
    .CLK(dco_clk),
    .D(_03422_),
    .Q( execution_unit_0.inst_dext_8_ ),
    .R(_03313_),
    .S(1'h1)
  );
  DFFSR _11290_ (
    .CLK(dco_clk),
    .D(_03423_),
    .Q( execution_unit_0.inst_dext_9_ ),
    .R(_03314_),
    .S(1'h1)
  );
  DFFSR _11291_ (
    .CLK(dco_clk),
    .D(_03424_),
    .Q( execution_unit_0.inst_dext_10_ ),
    .R(_03315_),
    .S(1'h1)
  );
  DFFSR _11292_ (
    .CLK(dco_clk),
    .D(_03425_),
    .Q( execution_unit_0.inst_dext_11_ ),
    .R(_03316_),
    .S(1'h1)
  );
  DFFSR _11293_ (
    .CLK(dco_clk),
    .D(_03426_),
    .Q( execution_unit_0.inst_dext_12_ ),
    .R(_03317_),
    .S(1'h1)
  );
  DFFSR _11294_ (
    .CLK(dco_clk),
    .D(_03427_),
    .Q( execution_unit_0.inst_dext_13_ ),
    .R(_03318_),
    .S(1'h1)
  );
  DFFSR _11295_ (
    .CLK(dco_clk),
    .D(_03428_),
    .Q( execution_unit_0.inst_dext_14_ ),
    .R(_03319_),
    .S(1'h1)
  );
  DFFSR _11296_ (
    .CLK(dco_clk),
    .D(_03429_),
    .Q( execution_unit_0.inst_dext_15_ ),
    .R(_03320_),
    .S(1'h1)
  );
  DFFSR _11297_ (
    .CLK(dco_clk),
    .D( frontend_0.fe_pmem_wait ),
    .Q( frontend_0.pmem_busy ),
    .R(_03321_),
    .S(1'h1)
  );
  DFFSR _11298_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_0_ ),
    .Q( dbg_0.UNUSED_pc_0_ ),
    .R(_03322_),
    .S(1'h1)
  );
  DFFSR _11299_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_1_ ),
    .Q( dbg_0.UNUSED_pc_1_ ),
    .R(_03323_),
    .S(1'h1)
  );
  DFFSR _11300_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_2_ ),
    .Q( dbg_0.UNUSED_pc_2_ ),
    .R(_03324_),
    .S(1'h1)
  );
  DFFSR _11301_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_3_ ),
    .Q( dbg_0.UNUSED_pc_3_ ),
    .R(_03325_),
    .S(1'h1)
  );
  DFFSR _11302_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_4_ ),
    .Q( dbg_0.UNUSED_pc_4_ ),
    .R(_03326_),
    .S(1'h1)
  );
  DFFSR _11303_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_5_ ),
    .Q( dbg_0.UNUSED_pc_5_ ),
    .R(_03327_),
    .S(1'h1)
  );
  DFFSR _11304_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_6_ ),
    .Q( dbg_0.UNUSED_pc_6_ ),
    .R(_03328_),
    .S(1'h1)
  );
  DFFSR _11305_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_7_ ),
    .Q( dbg_0.UNUSED_pc_7_ ),
    .R(_03329_),
    .S(1'h1)
  );
  DFFSR _11306_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_8_ ),
    .Q( dbg_0.UNUSED_pc_8_ ),
    .R(_03330_),
    .S(1'h1)
  );
  DFFSR _11307_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_9_ ),
    .Q( dbg_0.UNUSED_pc_9_ ),
    .R(_03331_),
    .S(1'h1)
  );
  DFFSR _11308_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_10_ ),
    .Q( dbg_0.UNUSED_pc_10_ ),
    .R(_03332_),
    .S(1'h1)
  );
  DFFSR _11309_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_11_ ),
    .Q( dbg_0.UNUSED_pc_11_ ),
    .R(_03333_),
    .S(1'h1)
  );
  DFFSR _11310_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_12_ ),
    .Q( dbg_0.UNUSED_pc_12_ ),
    .R(_03334_),
    .S(1'h1)
  );
  DFFSR _11311_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_13_ ),
    .Q( dbg_0.UNUSED_pc_13_ ),
    .R(_03335_),
    .S(1'h1)
  );
  DFFSR _11312_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_14_ ),
    .Q( dbg_0.UNUSED_pc_14_ ),
    .R(_03336_),
    .S(1'h1)
  );
  DFFSR _11313_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_15_ ),
    .Q( dbg_0.UNUSED_pc_15_ ),
    .R(_03337_),
    .S(1'h1)
  );
  DFFSR _11314_ (
    .CLK(dco_clk),
    .D(_03430_),
    .Q( execution_unit_0.inst_sext_0_ ),
    .R(_03338_),
    .S(1'h1)
  );
  DFFSR _11315_ (
    .CLK(dco_clk),
    .D(_03431_),
    .Q( execution_unit_0.inst_sext_1_ ),
    .R(_03339_),
    .S(1'h1)
  );
  DFFSR _11316_ (
    .CLK(dco_clk),
    .D(_03432_),
    .Q( execution_unit_0.inst_sext_2_ ),
    .R(_03340_),
    .S(1'h1)
  );
  DFFSR _11317_ (
    .CLK(dco_clk),
    .D(_03433_),
    .Q( execution_unit_0.inst_sext_3_ ),
    .R(_03341_),
    .S(1'h1)
  );
  DFFSR _11318_ (
    .CLK(dco_clk),
    .D(_03434_),
    .Q( execution_unit_0.inst_sext_4_ ),
    .R(_03342_),
    .S(1'h1)
  );
  DFFSR _11319_ (
    .CLK(dco_clk),
    .D(_03435_),
    .Q( execution_unit_0.inst_sext_5_ ),
    .R(_03343_),
    .S(1'h1)
  );
  DFFSR _11320_ (
    .CLK(dco_clk),
    .D(_03436_),
    .Q( execution_unit_0.inst_sext_6_ ),
    .R(_03344_),
    .S(1'h1)
  );
  DFFSR _11321_ (
    .CLK(dco_clk),
    .D(_03437_),
    .Q( execution_unit_0.inst_sext_7_ ),
    .R(_03345_),
    .S(1'h1)
  );
  DFFSR _11322_ (
    .CLK(dco_clk),
    .D(_03438_),
    .Q( execution_unit_0.inst_sext_8_ ),
    .R(_03346_),
    .S(1'h1)
  );
  DFFSR _11323_ (
    .CLK(dco_clk),
    .D(_03439_),
    .Q( execution_unit_0.inst_sext_9_ ),
    .R(_03347_),
    .S(1'h1)
  );
  DFFSR _11324_ (
    .CLK(dco_clk),
    .D(_03440_),
    .Q( execution_unit_0.inst_sext_10_ ),
    .R(_03348_),
    .S(1'h1)
  );
  DFFSR _11325_ (
    .CLK(dco_clk),
    .D(_03441_),
    .Q( execution_unit_0.inst_sext_11_ ),
    .R(_03349_),
    .S(1'h1)
  );
  DFFSR _11326_ (
    .CLK(dco_clk),
    .D(_03442_),
    .Q( execution_unit_0.inst_sext_12_ ),
    .R(_03350_),
    .S(1'h1)
  );
  DFFSR _11327_ (
    .CLK(dco_clk),
    .D(_03443_),
    .Q( execution_unit_0.inst_sext_13_ ),
    .R(_03351_),
    .S(1'h1)
  );
  DFFSR _11328_ (
    .CLK(dco_clk),
    .D(_03444_),
    .Q( execution_unit_0.inst_sext_14_ ),
    .R(_03352_),
    .S(1'h1)
  );
  DFFSR _11329_ (
    .CLK(dco_clk),
    .D(_03445_),
    .Q( execution_unit_0.inst_sext_15_ ),
    .R(_03353_),
    .S(1'h1)
  );
  DFFSR _11330_ (
    .CLK(dco_clk),
    .D(_03446_),
    .Q( execution_unit_0.inst_ad_0_ ),
    .R(_03354_),
    .S(1'h1)
  );
  DFFSR _11331_ (
    .CLK(dco_clk),
    .D(_03447_),
    .Q( execution_unit_0.UNUSED_inst_ad_idx ),
    .R(_03355_),
    .S(1'h1)
  );
  DFFSR _11332_ (
    .CLK(dco_clk),
    .D(_03448_),
    .Q( execution_unit_0.UNUSED_inst_ad_symb ),
    .R(_03356_),
    .S(1'h1)
  );
  DFFSR _11333_ (
    .CLK(dco_clk),
    .D(_03449_),
    .Q( execution_unit_0.inst_ad_6_ ),
    .R(_03357_),
    .S(1'h1)
  );
  DFFSR _11334_ (
    .CLK(dco_clk),
    .D(_03253_),
    .Q( dbg_0.cpu_stat_full_0_ ),
    .R(_03358_),
    .S(1'h1)
  );
  DFFSR _11335_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_0_ ),
    .Q( frontend_0.i_state_0_ ),
    .R(_03359_),
    .S(1'h1)
  );
  DFFSR _11336_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_1_ ),
    .Q( frontend_0.i_state_1_ ),
    .R(_03360_),
    .S(1'h1)
  );
  DFFSR _11337_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_2_ ),
    .Q( frontend_0.i_state_2_ ),
    .R(_03361_),
    .S(1'h1)
  );
  DFFSR _11338_ (
    .CLK(dco_clk),
    .D(_03450_),
    .Q( execution_unit_0.inst_irq_rst ),
    .R(1'h1),
    .S(_03362_)
  );
  DFFSR _11339_ (
    .CLK(dco_clk),
    .D(_03451_),
    .Q( frontend_0.irq_addr_1_ ),
    .R(1'h1),
    .S(_03363_)
  );
  DFFSR _11340_ (
    .CLK(dco_clk),
    .D(_03452_),
    .Q( frontend_0.irq_addr_2_ ),
    .R(1'h1),
    .S(_03364_)
  );
  DFFSR _11341_ (
    .CLK(dco_clk),
    .D(_03453_),
    .Q( frontend_0.irq_addr_3_ ),
    .R(1'h1),
    .S(_03365_)
  );
  DFFSR _11342_ (
    .CLK(dco_clk),
    .D(_03454_),
    .Q( frontend_0.irq_addr_4_ ),
    .R(1'h1),
    .S(_03366_)
  );
  INVX1 _11343_ (
    .A(pmem_dout_15_),
    .Y(_04257_)
  );
  INVX1 _11344_ (
    .A(pmem_dout_14_),
    .Y(_04258_)
  );
  INVX1 _11345_ (
    .A(pmem_dout_13_),
    .Y(_04259_)
  );
  INVX1 _11346_ (
    .A(pmem_dout_12_),
    .Y(_04260_)
  );
  INVX1 _11347_ (
    .A(pmem_dout_11_),
    .Y(_04261_)
  );
  INVX1 _11348_ (
    .A(pmem_dout_10_),
    .Y(_04262_)
  );
  INVX1 _11349_ (
    .A(pmem_dout_9_),
    .Y(_04263_)
  );
  INVX1 _11350_ (
    .A(pmem_dout_8_),
    .Y(_04264_)
  );
  INVX1 _11351_ (
    .A(pmem_dout_7_),
    .Y(_04265_)
  );
  INVX1 _11352_ (
    .A(pmem_dout_6_),
    .Y(_04266_)
  );
  INVX1 _11353_ (
    .A(pmem_dout_5_),
    .Y(_04267_)
  );
  INVX1 _11354_ (
    .A(pmem_dout_4_),
    .Y(_04268_)
  );
  INVX1 _11355_ (
    .A(pmem_dout_3_),
    .Y(_04269_)
  );
  INVX1 _11356_ (
    .A(pmem_dout_2_),
    .Y(_04270_)
  );
  INVX1 _11357_ (
    .A(pmem_dout_1_),
    .Y(_04271_)
  );
  INVX1 _11358_ (
    .A(pmem_dout_0_),
    .Y(_04272_)
  );
  INVX1 _11359_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_04273_)
  );
  INVX1 _11360_ (
    .A( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .Y(_04274_)
  );
  INVX1 _11361_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .Y(_04275_)
  );
  INVX1 _11362_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .Y(_04276_)
  );
  INVX1 _11363_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .Y(_04277_)
  );
  INVX1 _11364_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .Y(_04278_)
  );
  INVX1 _11365_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .Y(_04279_)
  );
  INVX1 _11366_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .Y(_04280_)
  );
  INVX1 _11367_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .Y(_04281_)
  );
  INVX1 _11368_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .Y(_04282_)
  );
  INVX1 _11369_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .Y(_04283_)
  );
  INVX1 _11370_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .Y(_04284_)
  );
  INVX1 _11371_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .Y(_04285_)
  );
  INVX1 _11372_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .Y(_04286_)
  );
  INVX1 _11373_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .Y(_04287_)
  );
  INVX1 _11374_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .Y(_04288_)
  );
  INVX1 _11375_ (
    .A( dbg_0.dbg_mem_addr_7_ ),
    .Y(_04289_)
  );
  INVX1 _11376_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .Y(_04290_)
  );
  INVX1 _11377_ (
    .A( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_04291_)
  );
  INVX1 _11378_ (
    .A( dbg_0.UNUSED_eu_mab_10_ ),
    .Y(_04292_)
  );
  INVX1 _11379_ (
    .A( dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_04293_)
  );
  INVX1 _11380_ (
    .A( dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_04294_)
  );
  INVX1 _11381_ (
    .A( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_04295_)
  );
  INVX1 _11382_ (
    .A( dbg_0.UNUSED_eu_mab_6_ ),
    .Y(_04296_)
  );
  INVX1 _11383_ (
    .A( dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_04297_)
  );
  INVX1 _11384_ (
    .A( dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_04298_)
  );
  INVX1 _11385_ (
    .A( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_04299_)
  );
  INVX1 _11386_ (
    .A( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_04300_)
  );
  INVX1 _11387_ (
    .A( dbg_0.UNUSED_eu_mab_1_ ),
    .Y(_04301_)
  );
  INVX1 _11388_ (
    .A( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_04302_)
  );
  INVX1 _11389_ (
    .A( dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_04303_)
  );
  INVX1 _11390_ (
    .A( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_04304_)
  );
  INVX1 _11391_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .Y(_04305_)
  );
  INVX1 _11392_ (
    .A(_06309_),
    .Y(_04306_)
  );
  INVX1 _11393_ (
    .A( execution_unit_0.mdb_out_0_ ),
    .Y(_04307_)
  );
  INVX1 _11394_ (
    .A(_06316_),
    .Y(_04308_)
  );
  INVX1 _11395_ (
    .A( execution_unit_0.mdb_out_1_ ),
    .Y(_04309_)
  );
  INVX1 _11396_ (
    .A(_06317_),
    .Y(_04310_)
  );
  INVX1 _11397_ (
    .A( execution_unit_0.mdb_out_2_ ),
    .Y(_04311_)
  );
  INVX1 _11398_ (
    .A(_06318_),
    .Y(_04312_)
  );
  INVX1 _11399_ (
    .A( execution_unit_0.mdb_out_3_ ),
    .Y(_04313_)
  );
  INVX1 _11400_ (
    .A(_06319_),
    .Y(_04314_)
  );
  INVX1 _11401_ (
    .A( execution_unit_0.mdb_out_4_ ),
    .Y(_04315_)
  );
  INVX1 _11402_ (
    .A(_06320_),
    .Y(_04316_)
  );
  INVX1 _11403_ (
    .A( execution_unit_0.mdb_out_5_ ),
    .Y(_04317_)
  );
  INVX1 _11404_ (
    .A(_06321_),
    .Y(_04318_)
  );
  INVX1 _11405_ (
    .A( execution_unit_0.mdb_out_6_ ),
    .Y(_04319_)
  );
  INVX1 _11406_ (
    .A(_06322_),
    .Y(_04320_)
  );
  INVX1 _11407_ (
    .A( execution_unit_0.mdb_out_7_ ),
    .Y(_04321_)
  );
  INVX1 _11408_ (
    .A(_06323_),
    .Y(_04322_)
  );
  INVX1 _11409_ (
    .A( execution_unit_0.mdb_out_8_ ),
    .Y(_04323_)
  );
  INVX1 _11410_ (
    .A(_06324_),
    .Y(_04324_)
  );
  INVX1 _11411_ (
    .A( execution_unit_0.mdb_out_9_ ),
    .Y(_04325_)
  );
  INVX1 _11412_ (
    .A(_06310_),
    .Y(_04326_)
  );
  INVX1 _11413_ (
    .A( execution_unit_0.mdb_out_10_ ),
    .Y(_04327_)
  );
  INVX1 _11414_ (
    .A(_06311_),
    .Y(_04328_)
  );
  INVX1 _11415_ (
    .A( execution_unit_0.mdb_out_11_ ),
    .Y(_04329_)
  );
  INVX1 _11416_ (
    .A(_06312_),
    .Y(_04330_)
  );
  INVX1 _11417_ (
    .A( execution_unit_0.mdb_out_12_ ),
    .Y(_04331_)
  );
  INVX1 _11418_ (
    .A(_06313_),
    .Y(_04332_)
  );
  INVX1 _11419_ (
    .A( execution_unit_0.mdb_out_13_ ),
    .Y(_04333_)
  );
  INVX1 _11420_ (
    .A(_06314_),
    .Y(_04334_)
  );
  INVX1 _11421_ (
    .A( execution_unit_0.mdb_out_14_ ),
    .Y(_04335_)
  );
  INVX1 _11422_ (
    .A(_06315_),
    .Y(_04336_)
  );
  INVX1 _11423_ (
    .A( execution_unit_0.mdb_out_15_ ),
    .Y(_04337_)
  );
  INVX1 _11424_ (
    .A(_06327_),
    .Y(_04202_)
  );
  NAND2X1 _11425_ (
    .A( frontend_0.mb_en ),
    .B( execution_unit_0.pc_nxt_15_ ),
    .Y(_04338_)
  );
  INVX1 _11426_ (
    .A(_04338_),
    .Y( mem_backbone_0.fe_pmem_en )
  );
  NAND3X1 _11427_ (
    .A( mem_backbone_0.fe_pmem_en_dly ),
    .B(_04273_),
    .C(_04338_),
    .Y(_04339_)
  );
  NOR2X1 _11428_ (
    .A( mem_backbone_0.fe_pmem_en_dly ),
    .B(_04338_),
    .Y(_04340_)
  );
  NAND2X1 _11429_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04273_),
    .Y(_04341_)
  );
  OAI21X1 _11430_ (
    .A(_04340_),
    .B(_04341_),
    .C(_04339_),
    .Y(_04256_)
  );
  MUX2X1 _11431_ (
    .A( mem_backbone_0.pmem_dout_bckup_15_ ),
    .B(pmem_dout_15_),
    .S(_04339_),
    .Y(_04342_)
  );
  INVX1 _11432_ (
    .A(_04342_),
    .Y(_04255_)
  );
  MUX2X1 _11433_ (
    .A( mem_backbone_0.pmem_dout_bckup_14_ ),
    .B(pmem_dout_14_),
    .S(_04339_),
    .Y(_04343_)
  );
  INVX1 _11434_ (
    .A(_04343_),
    .Y(_04254_)
  );
  MUX2X1 _11435_ (
    .A( mem_backbone_0.pmem_dout_bckup_13_ ),
    .B(pmem_dout_13_),
    .S(_04339_),
    .Y(_04344_)
  );
  INVX1 _11436_ (
    .A(_04344_),
    .Y(_04253_)
  );
  MUX2X1 _11437_ (
    .A( mem_backbone_0.pmem_dout_bckup_12_ ),
    .B(pmem_dout_12_),
    .S(_04339_),
    .Y(_04345_)
  );
  INVX1 _11438_ (
    .A(_04345_),
    .Y(_04252_)
  );
  MUX2X1 _11439_ (
    .A( mem_backbone_0.pmem_dout_bckup_11_ ),
    .B(pmem_dout_11_),
    .S(_04339_),
    .Y(_04346_)
  );
  INVX1 _11440_ (
    .A(_04346_),
    .Y(_04251_)
  );
  MUX2X1 _11441_ (
    .A( mem_backbone_0.pmem_dout_bckup_10_ ),
    .B(pmem_dout_10_),
    .S(_04339_),
    .Y(_04347_)
  );
  INVX1 _11442_ (
    .A(_04347_),
    .Y(_04250_)
  );
  MUX2X1 _11443_ (
    .A( mem_backbone_0.pmem_dout_bckup_9_ ),
    .B(pmem_dout_9_),
    .S(_04339_),
    .Y(_04348_)
  );
  INVX1 _11444_ (
    .A(_04348_),
    .Y(_04249_)
  );
  MUX2X1 _11445_ (
    .A( mem_backbone_0.pmem_dout_bckup_8_ ),
    .B(pmem_dout_8_),
    .S(_04339_),
    .Y(_04349_)
  );
  INVX1 _11446_ (
    .A(_04349_),
    .Y(_04248_)
  );
  MUX2X1 _11447_ (
    .A( mem_backbone_0.pmem_dout_bckup_7_ ),
    .B(pmem_dout_7_),
    .S(_04339_),
    .Y(_04350_)
  );
  INVX1 _11448_ (
    .A(_04350_),
    .Y(_04247_)
  );
  MUX2X1 _11449_ (
    .A( mem_backbone_0.pmem_dout_bckup_6_ ),
    .B(pmem_dout_6_),
    .S(_04339_),
    .Y(_04351_)
  );
  INVX1 _11450_ (
    .A(_04351_),
    .Y(_04246_)
  );
  MUX2X1 _11451_ (
    .A( mem_backbone_0.pmem_dout_bckup_5_ ),
    .B(pmem_dout_5_),
    .S(_04339_),
    .Y(_04352_)
  );
  INVX1 _11452_ (
    .A(_04352_),
    .Y(_04245_)
  );
  MUX2X1 _11453_ (
    .A( mem_backbone_0.pmem_dout_bckup_4_ ),
    .B(pmem_dout_4_),
    .S(_04339_),
    .Y(_04353_)
  );
  INVX1 _11454_ (
    .A(_04353_),
    .Y(_04244_)
  );
  MUX2X1 _11455_ (
    .A( mem_backbone_0.pmem_dout_bckup_3_ ),
    .B(pmem_dout_3_),
    .S(_04339_),
    .Y(_04354_)
  );
  INVX1 _11456_ (
    .A(_04354_),
    .Y(_04243_)
  );
  MUX2X1 _11457_ (
    .A( mem_backbone_0.pmem_dout_bckup_2_ ),
    .B(pmem_dout_2_),
    .S(_04339_),
    .Y(_04355_)
  );
  INVX1 _11458_ (
    .A(_04355_),
    .Y(_04242_)
  );
  MUX2X1 _11459_ (
    .A( mem_backbone_0.pmem_dout_bckup_1_ ),
    .B(pmem_dout_1_),
    .S(_04339_),
    .Y(_04356_)
  );
  INVX1 _11460_ (
    .A(_04356_),
    .Y(_04241_)
  );
  MUX2X1 _11461_ (
    .A( mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(pmem_dout_0_),
    .S(_04339_),
    .Y(_04357_)
  );
  INVX1 _11462_ (
    .A(_04357_),
    .Y(_04240_)
  );
  NAND2X1 _11463_ (
    .A( dbg_0.UNUSED_eu_mab_14_ ),
    .B( dbg_0.UNUSED_eu_mb_en ),
    .Y(_04358_)
  );
  NOR2X1 _11464_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B(_04358_),
    .Y(_04359_)
  );
  NAND3X1 _11465_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_04290_),
    .C( dbg_0.dbg_mem_en ),
    .Y(_04360_)
  );
  NOR2X1 _11466_ (
    .A(_04359_),
    .B(_04360_),
    .Y(_04361_)
  );
  MUX2X1 _11467_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .S(_04361_),
    .Y(_06246_)
  );
  MUX2X1 _11468_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .S(_04361_),
    .Y(_06247_)
  );
  MUX2X1 _11469_ (
    .A(_04283_),
    .B(_04301_),
    .S(_04361_),
    .Y(_06216_)
  );
  MUX2X1 _11470_ (
    .A(_04282_),
    .B(_04300_),
    .S(_04361_),
    .Y(_06220_)
  );
  MUX2X1 _11471_ (
    .A(_04285_),
    .B(_04303_),
    .S(_04361_),
    .Y(_06221_)
  );
  MUX2X1 _11472_ (
    .A(_04284_),
    .B(_04302_),
    .S(_04361_),
    .Y(_06222_)
  );
  MUX2X1 _11473_ (
    .A(_04287_),
    .B(_04297_),
    .S(_04361_),
    .Y(_06223_)
  );
  MUX2X1 _11474_ (
    .A(_04286_),
    .B(_04296_),
    .S(_04361_),
    .Y(_06224_)
  );
  MUX2X1 _11475_ (
    .A(_04289_),
    .B(_04299_),
    .S(_04361_),
    .Y(_06225_)
  );
  MUX2X1 _11476_ (
    .A(_04288_),
    .B(_04298_),
    .S(_04361_),
    .Y(_06226_)
  );
  MUX2X1 _11477_ (
    .A(_04279_),
    .B(_04293_),
    .S(_04361_),
    .Y(_06227_)
  );
  MUX2X1 _11478_ (
    .A(_04278_),
    .B(_04292_),
    .S(_04361_),
    .Y(_06228_)
  );
  MUX2X1 _11479_ (
    .A(_04281_),
    .B(_04295_),
    .S(_04361_),
    .Y(_06217_)
  );
  MUX2X1 _11480_ (
    .A(_04280_),
    .B(_04294_),
    .S(_04361_),
    .Y(_06218_)
  );
  MUX2X1 _11481_ (
    .A(_04276_),
    .B(_04291_),
    .S(_04361_),
    .Y(_06219_)
  );
  MUX2X1 _11482_ (
    .A(_04306_),
    .B(_04307_),
    .S(_04361_),
    .Y(_06230_)
  );
  MUX2X1 _11483_ (
    .A(_04308_),
    .B(_04309_),
    .S(_04361_),
    .Y(_06237_)
  );
  MUX2X1 _11484_ (
    .A(_04310_),
    .B(_04311_),
    .S(_04361_),
    .Y(_06238_)
  );
  MUX2X1 _11485_ (
    .A(_04312_),
    .B(_04313_),
    .S(_04361_),
    .Y(_06239_)
  );
  MUX2X1 _11486_ (
    .A(_04314_),
    .B(_04315_),
    .S(_04361_),
    .Y(_06240_)
  );
  MUX2X1 _11487_ (
    .A(_04316_),
    .B(_04317_),
    .S(_04361_),
    .Y(_06241_)
  );
  MUX2X1 _11488_ (
    .A(_04318_),
    .B(_04319_),
    .S(_04361_),
    .Y(_06242_)
  );
  MUX2X1 _11489_ (
    .A(_04320_),
    .B(_04321_),
    .S(_04361_),
    .Y(_06243_)
  );
  MUX2X1 _11490_ (
    .A(_04322_),
    .B(_04323_),
    .S(_04361_),
    .Y(_06244_)
  );
  MUX2X1 _11491_ (
    .A(_04324_),
    .B(_04325_),
    .S(_04361_),
    .Y(_06245_)
  );
  MUX2X1 _11492_ (
    .A(_04326_),
    .B(_04327_),
    .S(_04361_),
    .Y(_06231_)
  );
  MUX2X1 _11493_ (
    .A(_04328_),
    .B(_04329_),
    .S(_04361_),
    .Y(_06232_)
  );
  MUX2X1 _11494_ (
    .A(_04330_),
    .B(_04331_),
    .S(_04361_),
    .Y(_06233_)
  );
  MUX2X1 _11495_ (
    .A(_04332_),
    .B(_04333_),
    .S(_04361_),
    .Y(_06234_)
  );
  MUX2X1 _11496_ (
    .A(_04334_),
    .B(_04335_),
    .S(_04361_),
    .Y(_06235_)
  );
  MUX2X1 _11497_ (
    .A(_04336_),
    .B(_04337_),
    .S(_04361_),
    .Y(_06236_)
  );
  OR2X1 _11498_ (
    .A( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_04362_)
  );
  NAND2X1 _11499_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B( dbg_0.UNUSED_eu_mb_en ),
    .Y(_04363_)
  );
  NOR2X1 _11500_ (
    .A(_04362_),
    .B(_04363_),
    .Y( mem_backbone_0.eu_pmem_en )
  );
  OAI21X1 _11501_ (
    .A(_04362_),
    .B(_04363_),
    .C(_04338_),
    .Y(_04364_)
  );
  NAND2X1 _11502_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B( dbg_0.dbg_mem_en ),
    .Y(_04365_)
  );
  NOR2X1 _11503_ (
    .A(_04364_),
    .B(_04365_),
    .Y( mem_backbone_0.ext_pmem_en )
  );
  NAND2X1 _11504_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_06325_)
  );
  NAND2X1 _11505_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_06326_)
  );
  MUX2X1 _11506_ (
    .A( dbg_0.UNUSED_eu_mab_1_ ),
    .B( execution_unit_0.pc_nxt_1_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04366_)
  );
  MUX2X1 _11507_ (
    .A(_04283_),
    .B(_04366_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06294_)
  );
  MUX2X1 _11508_ (
    .A( dbg_0.UNUSED_eu_mab_2_ ),
    .B( execution_unit_0.pc_nxt_2_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04367_)
  );
  MUX2X1 _11509_ (
    .A(_04282_),
    .B(_04367_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06299_)
  );
  MUX2X1 _11510_ (
    .A( dbg_0.UNUSED_eu_mab_3_ ),
    .B( execution_unit_0.pc_nxt_3_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04368_)
  );
  MUX2X1 _11511_ (
    .A(_04285_),
    .B(_04368_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06300_)
  );
  MUX2X1 _11512_ (
    .A( dbg_0.UNUSED_eu_mab_4_ ),
    .B( execution_unit_0.pc_nxt_4_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04369_)
  );
  MUX2X1 _11513_ (
    .A(_04284_),
    .B(_04369_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06301_)
  );
  MUX2X1 _11514_ (
    .A( dbg_0.UNUSED_eu_mab_5_ ),
    .B( execution_unit_0.pc_nxt_5_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04370_)
  );
  MUX2X1 _11515_ (
    .A(_04287_),
    .B(_04370_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06302_)
  );
  MUX2X1 _11516_ (
    .A( dbg_0.UNUSED_eu_mab_6_ ),
    .B( execution_unit_0.pc_nxt_6_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04371_)
  );
  MUX2X1 _11517_ (
    .A(_04286_),
    .B(_04371_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06303_)
  );
  MUX2X1 _11518_ (
    .A( dbg_0.UNUSED_eu_mab_7_ ),
    .B( execution_unit_0.pc_nxt_7_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04372_)
  );
  MUX2X1 _11519_ (
    .A(_04289_),
    .B(_04372_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06304_)
  );
  MUX2X1 _11520_ (
    .A( dbg_0.UNUSED_eu_mab_8_ ),
    .B( execution_unit_0.pc_nxt_8_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04373_)
  );
  MUX2X1 _11521_ (
    .A(_04288_),
    .B(_04373_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06305_)
  );
  MUX2X1 _11522_ (
    .A( dbg_0.UNUSED_eu_mab_9_ ),
    .B( execution_unit_0.pc_nxt_9_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04374_)
  );
  MUX2X1 _11523_ (
    .A(_04279_),
    .B(_04374_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06306_)
  );
  MUX2X1 _11524_ (
    .A( dbg_0.UNUSED_eu_mab_10_ ),
    .B( execution_unit_0.pc_nxt_10_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04375_)
  );
  MUX2X1 _11525_ (
    .A(_04278_),
    .B(_04375_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06307_)
  );
  MUX2X1 _11526_ (
    .A( dbg_0.UNUSED_eu_mab_11_ ),
    .B( execution_unit_0.pc_nxt_11_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04376_)
  );
  MUX2X1 _11527_ (
    .A(_04281_),
    .B(_04376_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06295_)
  );
  MUX2X1 _11528_ (
    .A( dbg_0.UNUSED_eu_mab_12_ ),
    .B( execution_unit_0.pc_nxt_12_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04377_)
  );
  MUX2X1 _11529_ (
    .A(_04280_),
    .B(_04377_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06296_)
  );
  MUX2X1 _11530_ (
    .A( dbg_0.UNUSED_eu_mab_13_ ),
    .B( execution_unit_0.pc_nxt_13_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04378_)
  );
  MUX2X1 _11531_ (
    .A(_04276_),
    .B(_04378_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06297_)
  );
  MUX2X1 _11532_ (
    .A( dbg_0.UNUSED_eu_mab_14_ ),
    .B( execution_unit_0.pc_nxt_14_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_04379_)
  );
  MUX2X1 _11533_ (
    .A(_04277_),
    .B(_04379_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_06298_)
  );
  NOR2X1 _11534_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_04380_)
  );
  NAND2X1 _11535_ (
    .A( dbg_0.UNUSED_eu_mb_en ),
    .B(_04380_),
    .Y(_04381_)
  );
  INVX1 _11536_ (
    .A(_04381_),
    .Y( mem_backbone_0.eu_per_en )
  );
  NAND3X1 _11537_ (
    .A(_04277_),
    .B(_04290_),
    .C( dbg_0.dbg_mem_en ),
    .Y(_04382_)
  );
  NOR2X1 _11538_ (
    .A( mem_backbone_0.eu_per_en ),
    .B(_04382_),
    .Y( mem_backbone_0.ext_per_en )
  );
  MUX2X1 _11539_ (
    .A(_04275_),
    .B(_04274_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06292_)
  );
  MUX2X1 _11540_ (
    .A(_04305_),
    .B(_04304_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06293_)
  );
  MUX2X1 _11541_ (
    .A(_04283_),
    .B(_04301_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06262_)
  );
  MUX2X1 _11542_ (
    .A(_04282_),
    .B(_04300_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06266_)
  );
  MUX2X1 _11543_ (
    .A(_04285_),
    .B(_04303_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06267_)
  );
  MUX2X1 _11544_ (
    .A(_04284_),
    .B(_04302_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06268_)
  );
  MUX2X1 _11545_ (
    .A(_04287_),
    .B(_04297_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06269_)
  );
  MUX2X1 _11546_ (
    .A(_04286_),
    .B(_04296_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06270_)
  );
  MUX2X1 _11547_ (
    .A(_04289_),
    .B(_04299_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06271_)
  );
  MUX2X1 _11548_ (
    .A(_04288_),
    .B(_04298_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06272_)
  );
  MUX2X1 _11549_ (
    .A(_04279_),
    .B(_04293_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06273_)
  );
  MUX2X1 _11550_ (
    .A(_04278_),
    .B(_04292_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06274_)
  );
  MUX2X1 _11551_ (
    .A(_04281_),
    .B(_04295_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06263_)
  );
  MUX2X1 _11552_ (
    .A(_04280_),
    .B(_04294_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06264_)
  );
  MUX2X1 _11553_ (
    .A(_04276_),
    .B(_04291_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06265_)
  );
  MUX2X1 _11554_ (
    .A(_04306_),
    .B(_04307_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06275_)
  );
  MUX2X1 _11555_ (
    .A(_04308_),
    .B(_04309_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06282_)
  );
  MUX2X1 _11556_ (
    .A(_04310_),
    .B(_04311_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06283_)
  );
  MUX2X1 _11557_ (
    .A(_04312_),
    .B(_04313_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06284_)
  );
  MUX2X1 _11558_ (
    .A(_04314_),
    .B(_04315_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06285_)
  );
  MUX2X1 _11559_ (
    .A(_04316_),
    .B(_04317_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06286_)
  );
  MUX2X1 _11560_ (
    .A(_04318_),
    .B(_04319_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06287_)
  );
  MUX2X1 _11561_ (
    .A(_04320_),
    .B(_04321_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06288_)
  );
  MUX2X1 _11562_ (
    .A(_04322_),
    .B(_04323_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06289_)
  );
  MUX2X1 _11563_ (
    .A(_04324_),
    .B(_04325_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06290_)
  );
  MUX2X1 _11564_ (
    .A(_04326_),
    .B(_04327_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06276_)
  );
  MUX2X1 _11565_ (
    .A(_04328_),
    .B(_04329_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06277_)
  );
  MUX2X1 _11566_ (
    .A(_04330_),
    .B(_04331_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06278_)
  );
  MUX2X1 _11567_ (
    .A(_04332_),
    .B(_04333_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06279_)
  );
  MUX2X1 _11568_ (
    .A(_04334_),
    .B(_04335_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06280_)
  );
  MUX2X1 _11569_ (
    .A(_04336_),
    .B(_04337_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_06281_)
  );
  NAND2X1 _11570_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_0_ ),
    .Y(_04383_)
  );
  OAI21X1 _11571_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04272_),
    .C(_04383_),
    .Y( dbg_0.fe_mdb_in_0_ )
  );
  NAND2X1 _11572_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_1_ ),
    .Y(_04384_)
  );
  OAI21X1 _11573_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04271_),
    .C(_04384_),
    .Y( dbg_0.fe_mdb_in_1_ )
  );
  NAND2X1 _11574_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_2_ ),
    .Y(_04385_)
  );
  OAI21X1 _11575_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04270_),
    .C(_04385_),
    .Y( dbg_0.fe_mdb_in_2_ )
  );
  NAND2X1 _11576_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_3_ ),
    .Y(_04386_)
  );
  OAI21X1 _11577_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04269_),
    .C(_04386_),
    .Y( dbg_0.fe_mdb_in_3_ )
  );
  NAND2X1 _11578_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_4_ ),
    .Y(_04387_)
  );
  OAI21X1 _11579_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04268_),
    .C(_04387_),
    .Y( dbg_0.fe_mdb_in_4_ )
  );
  NAND2X1 _11580_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_5_ ),
    .Y(_04388_)
  );
  OAI21X1 _11581_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04267_),
    .C(_04388_),
    .Y( dbg_0.fe_mdb_in_5_ )
  );
  NAND2X1 _11582_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_6_ ),
    .Y(_04389_)
  );
  OAI21X1 _11583_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04266_),
    .C(_04389_),
    .Y( dbg_0.fe_mdb_in_6_ )
  );
  NAND2X1 _11584_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_7_ ),
    .Y(_04390_)
  );
  OAI21X1 _11585_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04265_),
    .C(_04390_),
    .Y( dbg_0.fe_mdb_in_7_ )
  );
  NAND2X1 _11586_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_8_ ),
    .Y(_04391_)
  );
  OAI21X1 _11587_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04264_),
    .C(_04391_),
    .Y( dbg_0.fe_mdb_in_8_ )
  );
  NAND2X1 _11588_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_9_ ),
    .Y(_04392_)
  );
  OAI21X1 _11589_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04263_),
    .C(_04392_),
    .Y( dbg_0.fe_mdb_in_9_ )
  );
  NAND2X1 _11590_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_10_ ),
    .Y(_04393_)
  );
  OAI21X1 _11591_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04262_),
    .C(_04393_),
    .Y( dbg_0.fe_mdb_in_10_ )
  );
  NAND2X1 _11592_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_11_ ),
    .Y(_04394_)
  );
  OAI21X1 _11593_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04261_),
    .C(_04394_),
    .Y( dbg_0.fe_mdb_in_11_ )
  );
  NAND2X1 _11594_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_12_ ),
    .Y(_04395_)
  );
  OAI21X1 _11595_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04260_),
    .C(_04395_),
    .Y( dbg_0.fe_mdb_in_12_ )
  );
  NAND2X1 _11596_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_13_ ),
    .Y(_04396_)
  );
  OAI21X1 _11597_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04259_),
    .C(_04396_),
    .Y( dbg_0.fe_mdb_in_13_ )
  );
  NAND2X1 _11598_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_14_ ),
    .Y(_04397_)
  );
  OAI21X1 _11599_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04258_),
    .C(_04397_),
    .Y( dbg_0.fe_mdb_in_14_ )
  );
  NAND2X1 _11600_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_15_ ),
    .Y(_04398_)
  );
  OAI21X1 _11601_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04257_),
    .C(_04398_),
    .Y( dbg_0.fe_mdb_in_15_ )
  );
  MUX2X1 _11602_ (
    .A( mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04399_)
  );
  NAND2X1 _11603_ (
    .A(pmem_dout_0_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04400_)
  );
  OAI21X1 _11604_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04399_),
    .C(_04400_),
    .Y( execution_unit_0.mdb_in_0_ )
  );
  MUX2X1 _11605_ (
    .A( mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04401_)
  );
  NAND2X1 _11606_ (
    .A(pmem_dout_1_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04402_)
  );
  OAI21X1 _11607_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04401_),
    .C(_04402_),
    .Y( execution_unit_0.mdb_in_1_ )
  );
  MUX2X1 _11608_ (
    .A( mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04403_)
  );
  NAND2X1 _11609_ (
    .A(pmem_dout_2_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04404_)
  );
  OAI21X1 _11610_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04403_),
    .C(_04404_),
    .Y( execution_unit_0.mdb_in_2_ )
  );
  MUX2X1 _11611_ (
    .A( mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04405_)
  );
  NAND2X1 _11612_ (
    .A(pmem_dout_3_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04406_)
  );
  OAI21X1 _11613_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04405_),
    .C(_04406_),
    .Y( execution_unit_0.mdb_in_3_ )
  );
  MUX2X1 _11614_ (
    .A( mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04407_)
  );
  NAND2X1 _11615_ (
    .A(pmem_dout_4_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04408_)
  );
  OAI21X1 _11616_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04407_),
    .C(_04408_),
    .Y( execution_unit_0.mdb_in_4_ )
  );
  MUX2X1 _11617_ (
    .A( mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04409_)
  );
  NAND2X1 _11618_ (
    .A(pmem_dout_5_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04410_)
  );
  OAI21X1 _11619_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04409_),
    .C(_04410_),
    .Y( execution_unit_0.mdb_in_5_ )
  );
  MUX2X1 _11620_ (
    .A( mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04411_)
  );
  NAND2X1 _11621_ (
    .A(pmem_dout_6_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04412_)
  );
  OAI21X1 _11622_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04411_),
    .C(_04412_),
    .Y( execution_unit_0.mdb_in_6_ )
  );
  MUX2X1 _11623_ (
    .A( mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04413_)
  );
  NAND2X1 _11624_ (
    .A(pmem_dout_7_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04414_)
  );
  OAI21X1 _11625_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04413_),
    .C(_04414_),
    .Y( execution_unit_0.mdb_in_7_ )
  );
  MUX2X1 _11626_ (
    .A( mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04415_)
  );
  NAND2X1 _11627_ (
    .A(pmem_dout_8_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04416_)
  );
  OAI21X1 _11628_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04415_),
    .C(_04416_),
    .Y( execution_unit_0.mdb_in_8_ )
  );
  MUX2X1 _11629_ (
    .A( mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04417_)
  );
  NAND2X1 _11630_ (
    .A(pmem_dout_9_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04418_)
  );
  OAI21X1 _11631_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04417_),
    .C(_04418_),
    .Y( execution_unit_0.mdb_in_9_ )
  );
  MUX2X1 _11632_ (
    .A( mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04419_)
  );
  NAND2X1 _11633_ (
    .A(pmem_dout_10_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04420_)
  );
  OAI21X1 _11634_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04419_),
    .C(_04420_),
    .Y( execution_unit_0.mdb_in_10_ )
  );
  MUX2X1 _11635_ (
    .A( mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04421_)
  );
  NAND2X1 _11636_ (
    .A(pmem_dout_11_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04422_)
  );
  OAI21X1 _11637_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04421_),
    .C(_04422_),
    .Y( execution_unit_0.mdb_in_11_ )
  );
  MUX2X1 _11638_ (
    .A( mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04423_)
  );
  NAND2X1 _11639_ (
    .A(pmem_dout_12_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04424_)
  );
  OAI21X1 _11640_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04423_),
    .C(_04424_),
    .Y( execution_unit_0.mdb_in_12_ )
  );
  MUX2X1 _11641_ (
    .A( mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04425_)
  );
  NAND2X1 _11642_ (
    .A(pmem_dout_13_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04426_)
  );
  OAI21X1 _11643_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04425_),
    .C(_04426_),
    .Y( execution_unit_0.mdb_in_13_ )
  );
  MUX2X1 _11644_ (
    .A( mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04427_)
  );
  NAND2X1 _11645_ (
    .A(pmem_dout_14_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04428_)
  );
  OAI21X1 _11646_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04427_),
    .C(_04428_),
    .Y( execution_unit_0.mdb_in_14_ )
  );
  MUX2X1 _11647_ (
    .A( mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04429_)
  );
  NAND2X1 _11648_ (
    .A(pmem_dout_15_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04430_)
  );
  OAI21X1 _11649_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04429_),
    .C(_04430_),
    .Y( execution_unit_0.mdb_in_15_ )
  );
  MUX2X1 _11650_ (
    .A( mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04431_)
  );
  NAND2X1 _11651_ (
    .A(pmem_dout_0_),
    .B(_04201_),
    .Y(_04432_)
  );
  OAI21X1 _11652_ (
    .A(_04201_),
    .B(_04431_),
    .C(_04432_),
    .Y( dbg_0.dbg_mem_din_0_ )
  );
  MUX2X1 _11653_ (
    .A( mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04433_)
  );
  NAND2X1 _11654_ (
    .A(pmem_dout_1_),
    .B(_04201_),
    .Y(_04434_)
  );
  OAI21X1 _11655_ (
    .A(_04201_),
    .B(_04433_),
    .C(_04434_),
    .Y( dbg_0.dbg_mem_din_1_ )
  );
  MUX2X1 _11656_ (
    .A( mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04435_)
  );
  NAND2X1 _11657_ (
    .A(pmem_dout_2_),
    .B(_04201_),
    .Y(_04436_)
  );
  OAI21X1 _11658_ (
    .A(_04201_),
    .B(_04435_),
    .C(_04436_),
    .Y( dbg_0.dbg_mem_din_2_ )
  );
  MUX2X1 _11659_ (
    .A( mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04437_)
  );
  NAND2X1 _11660_ (
    .A(pmem_dout_3_),
    .B(_04201_),
    .Y(_04438_)
  );
  OAI21X1 _11661_ (
    .A(_04201_),
    .B(_04437_),
    .C(_04438_),
    .Y( dbg_0.dbg_mem_din_3_ )
  );
  MUX2X1 _11662_ (
    .A( mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04439_)
  );
  NAND2X1 _11663_ (
    .A(pmem_dout_4_),
    .B(_04201_),
    .Y(_04440_)
  );
  OAI21X1 _11664_ (
    .A(_04201_),
    .B(_04439_),
    .C(_04440_),
    .Y( dbg_0.dbg_mem_din_4_ )
  );
  MUX2X1 _11665_ (
    .A( mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04441_)
  );
  NAND2X1 _11666_ (
    .A(pmem_dout_5_),
    .B(_04201_),
    .Y(_04442_)
  );
  OAI21X1 _11667_ (
    .A(_04201_),
    .B(_04441_),
    .C(_04442_),
    .Y( dbg_0.dbg_mem_din_5_ )
  );
  MUX2X1 _11668_ (
    .A( mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04443_)
  );
  NAND2X1 _11669_ (
    .A(pmem_dout_6_),
    .B(_04201_),
    .Y(_04444_)
  );
  OAI21X1 _11670_ (
    .A(_04201_),
    .B(_04443_),
    .C(_04444_),
    .Y( dbg_0.dbg_mem_din_6_ )
  );
  MUX2X1 _11671_ (
    .A( mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04445_)
  );
  NAND2X1 _11672_ (
    .A(pmem_dout_7_),
    .B(_04201_),
    .Y(_04446_)
  );
  OAI21X1 _11673_ (
    .A(_04201_),
    .B(_04445_),
    .C(_04446_),
    .Y( dbg_0.dbg_mem_din_7_ )
  );
  MUX2X1 _11674_ (
    .A( mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04447_)
  );
  NAND2X1 _11675_ (
    .A(pmem_dout_8_),
    .B(_04201_),
    .Y(_04448_)
  );
  OAI21X1 _11676_ (
    .A(_04201_),
    .B(_04447_),
    .C(_04448_),
    .Y( dbg_0.dbg_mem_din_8_ )
  );
  MUX2X1 _11677_ (
    .A( mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04449_)
  );
  NAND2X1 _11678_ (
    .A(pmem_dout_9_),
    .B(_04201_),
    .Y(_04450_)
  );
  OAI21X1 _11679_ (
    .A(_04201_),
    .B(_04449_),
    .C(_04450_),
    .Y( dbg_0.dbg_mem_din_9_ )
  );
  MUX2X1 _11680_ (
    .A( mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04451_)
  );
  NAND2X1 _11681_ (
    .A(pmem_dout_10_),
    .B(_04201_),
    .Y(_04452_)
  );
  OAI21X1 _11682_ (
    .A(_04201_),
    .B(_04451_),
    .C(_04452_),
    .Y( dbg_0.dbg_mem_din_10_ )
  );
  MUX2X1 _11683_ (
    .A( mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04453_)
  );
  NAND2X1 _11684_ (
    .A(pmem_dout_11_),
    .B(_04201_),
    .Y(_04454_)
  );
  OAI21X1 _11685_ (
    .A(_04201_),
    .B(_04453_),
    .C(_04454_),
    .Y( dbg_0.dbg_mem_din_11_ )
  );
  MUX2X1 _11686_ (
    .A( mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04455_)
  );
  NAND2X1 _11687_ (
    .A(pmem_dout_12_),
    .B(_04201_),
    .Y(_04456_)
  );
  OAI21X1 _11688_ (
    .A(_04201_),
    .B(_04455_),
    .C(_04456_),
    .Y( dbg_0.dbg_mem_din_12_ )
  );
  MUX2X1 _11689_ (
    .A( mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04457_)
  );
  NAND2X1 _11690_ (
    .A(pmem_dout_13_),
    .B(_04201_),
    .Y(_04458_)
  );
  OAI21X1 _11691_ (
    .A(_04201_),
    .B(_04457_),
    .C(_04458_),
    .Y( dbg_0.dbg_mem_din_13_ )
  );
  MUX2X1 _11692_ (
    .A( mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04459_)
  );
  NAND2X1 _11693_ (
    .A(pmem_dout_14_),
    .B(_04201_),
    .Y(_04460_)
  );
  OAI21X1 _11694_ (
    .A(_04201_),
    .B(_04459_),
    .C(_04460_),
    .Y( dbg_0.dbg_mem_din_14_ )
  );
  MUX2X1 _11695_ (
    .A( mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_04461_)
  );
  NAND2X1 _11696_ (
    .A(pmem_dout_15_),
    .B(_04201_),
    .Y(_04462_)
  );
  OAI21X1 _11697_ (
    .A(_04201_),
    .B(_04461_),
    .C(_04462_),
    .Y( dbg_0.dbg_mem_din_15_ )
  );
  OAI21X1 _11698_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B(_04358_),
    .C(_04360_),
    .Y(_04463_)
  );
  INVX1 _11699_ (
    .A(_04463_),
    .Y(_06229_)
  );
  NOR2X1 _11700_ (
    .A(_04364_),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_06308_)
  );
  AND2X1 _11701_ (
    .A( mem_backbone_0.fe_pmem_en ),
    .B( mem_backbone_0.eu_pmem_en ),
    .Y( frontend_0.fe_pmem_wait )
  );
  NAND2X1 _11702_ (
    .A(_04381_),
    .B(_04382_),
    .Y(_06291_)
  );
  INVX1 _11703_ (
    .A(_06327_),
    .Y(_04203_)
  );
  INVX1 _11704_ (
    .A(_06327_),
    .Y(_04204_)
  );
  INVX1 _11705_ (
    .A(_06327_),
    .Y(_04205_)
  );
  INVX1 _11706_ (
    .A(_06327_),
    .Y(_04206_)
  );
  INVX1 _11707_ (
    .A(_06327_),
    .Y(_04207_)
  );
  INVX1 _11708_ (
    .A(_06327_),
    .Y(_04208_)
  );
  INVX1 _11709_ (
    .A(_06327_),
    .Y(_04209_)
  );
  INVX1 _11710_ (
    .A(_06327_),
    .Y(_04210_)
  );
  INVX1 _11711_ (
    .A(_06327_),
    .Y(_04211_)
  );
  INVX1 _11712_ (
    .A(_06327_),
    .Y(_04212_)
  );
  INVX1 _11713_ (
    .A(_06327_),
    .Y(_04213_)
  );
  INVX1 _11714_ (
    .A(_06327_),
    .Y(_04214_)
  );
  INVX1 _11715_ (
    .A(_06327_),
    .Y(_04215_)
  );
  INVX1 _11716_ (
    .A(_06327_),
    .Y(_04216_)
  );
  INVX1 _11717_ (
    .A(_06327_),
    .Y(_04217_)
  );
  INVX1 _11718_ (
    .A(_06327_),
    .Y(_04218_)
  );
  INVX1 _11719_ (
    .A(_06327_),
    .Y(_04219_)
  );
  INVX1 _11720_ (
    .A(_06327_),
    .Y(_04220_)
  );
  INVX1 _11721_ (
    .A(_06327_),
    .Y(_04221_)
  );
  INVX1 _11722_ (
    .A(_06327_),
    .Y(_04222_)
  );
  INVX1 _11723_ (
    .A(_06327_),
    .Y(_04223_)
  );
  INVX1 _11724_ (
    .A(_06327_),
    .Y(_04224_)
  );
  INVX1 _11725_ (
    .A(_06327_),
    .Y(_04225_)
  );
  INVX1 _11726_ (
    .A(_06327_),
    .Y(_04226_)
  );
  INVX1 _11727_ (
    .A(_06327_),
    .Y(_04227_)
  );
  INVX1 _11728_ (
    .A(_06327_),
    .Y(_04228_)
  );
  INVX1 _11729_ (
    .A(_06327_),
    .Y(_04229_)
  );
  INVX1 _11730_ (
    .A(_06327_),
    .Y(_04230_)
  );
  INVX1 _11731_ (
    .A(_06327_),
    .Y(_04231_)
  );
  INVX1 _11732_ (
    .A(_06327_),
    .Y(_04232_)
  );
  INVX1 _11733_ (
    .A(_06327_),
    .Y(_04233_)
  );
  INVX1 _11734_ (
    .A(_06327_),
    .Y(_04234_)
  );
  INVX1 _11735_ (
    .A(_06327_),
    .Y(_04235_)
  );
  INVX1 _11736_ (
    .A(_06327_),
    .Y(_04236_)
  );
  INVX1 _11737_ (
    .A(_06327_),
    .Y(_04237_)
  );
  INVX1 _11738_ (
    .A(_06327_),
    .Y(_04238_)
  );
  INVX1 _11739_ (
    .A(_06327_),
    .Y(_04239_)
  );
  DFFSR _11740_ (
    .CLK(dco_clk),
    .D(_04240_),
    .Q( mem_backbone_0.pmem_dout_bckup_0_ ),
    .R(_04202_),
    .S(1'h1)
  );
  DFFSR _11741_ (
    .CLK(dco_clk),
    .D(_04241_),
    .Q( mem_backbone_0.pmem_dout_bckup_1_ ),
    .R(_04203_),
    .S(1'h1)
  );
  DFFSR _11742_ (
    .CLK(dco_clk),
    .D(_04242_),
    .Q( mem_backbone_0.pmem_dout_bckup_2_ ),
    .R(_04204_),
    .S(1'h1)
  );
  DFFSR _11743_ (
    .CLK(dco_clk),
    .D(_04243_),
    .Q( mem_backbone_0.pmem_dout_bckup_3_ ),
    .R(_04205_),
    .S(1'h1)
  );
  DFFSR _11744_ (
    .CLK(dco_clk),
    .D(_04244_),
    .Q( mem_backbone_0.pmem_dout_bckup_4_ ),
    .R(_04206_),
    .S(1'h1)
  );
  DFFSR _11745_ (
    .CLK(dco_clk),
    .D(_04245_),
    .Q( mem_backbone_0.pmem_dout_bckup_5_ ),
    .R(_04207_),
    .S(1'h1)
  );
  DFFSR _11746_ (
    .CLK(dco_clk),
    .D(_04246_),
    .Q( mem_backbone_0.pmem_dout_bckup_6_ ),
    .R(_04208_),
    .S(1'h1)
  );
  DFFSR _11747_ (
    .CLK(dco_clk),
    .D(_04247_),
    .Q( mem_backbone_0.pmem_dout_bckup_7_ ),
    .R(_04209_),
    .S(1'h1)
  );
  DFFSR _11748_ (
    .CLK(dco_clk),
    .D(_04248_),
    .Q( mem_backbone_0.pmem_dout_bckup_8_ ),
    .R(_04210_),
    .S(1'h1)
  );
  DFFSR _11749_ (
    .CLK(dco_clk),
    .D(_04249_),
    .Q( mem_backbone_0.pmem_dout_bckup_9_ ),
    .R(_04211_),
    .S(1'h1)
  );
  DFFSR _11750_ (
    .CLK(dco_clk),
    .D(_04250_),
    .Q( mem_backbone_0.pmem_dout_bckup_10_ ),
    .R(_04212_),
    .S(1'h1)
  );
  DFFSR _11751_ (
    .CLK(dco_clk),
    .D(_04251_),
    .Q( mem_backbone_0.pmem_dout_bckup_11_ ),
    .R(_04213_),
    .S(1'h1)
  );
  DFFSR _11752_ (
    .CLK(dco_clk),
    .D(_04252_),
    .Q( mem_backbone_0.pmem_dout_bckup_12_ ),
    .R(_04214_),
    .S(1'h1)
  );
  DFFSR _11753_ (
    .CLK(dco_clk),
    .D(_04253_),
    .Q( mem_backbone_0.pmem_dout_bckup_13_ ),
    .R(_04215_),
    .S(1'h1)
  );
  DFFSR _11754_ (
    .CLK(dco_clk),
    .D(_04254_),
    .Q( mem_backbone_0.pmem_dout_bckup_14_ ),
    .R(_04216_),
    .S(1'h1)
  );
  DFFSR _11755_ (
    .CLK(dco_clk),
    .D(_04255_),
    .Q( mem_backbone_0.pmem_dout_bckup_15_ ),
    .R(_04217_),
    .S(1'h1)
  );
  DFFSR _11756_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.ext_per_en ),
    .Q( mem_backbone_0.ext_mem_din_sel ),
    .R(_04218_),
    .S(1'h1)
  );
  DFFSR _11757_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.ext_pmem_en ),
    .Q(_04201_),
    .R(_04219_),
    .S(1'h1)
  );
  DFFSR _11758_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.eu_per_en ),
    .Q( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .R(_04220_),
    .S(1'h1)
  );
  DFFSR _11759_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.eu_pmem_en ),
    .Q( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .R(_04221_),
    .S(1'h1)
  );
  DFFSR _11760_ (
    .CLK(dco_clk),
    .D(_04256_),
    .Q( mem_backbone_0.pmem_dout_bckup_sel ),
    .R(_04222_),
    .S(1'h1)
  );
  DFFSR _11761_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.fe_pmem_en ),
    .Q( mem_backbone_0.fe_pmem_en_dly ),
    .R(_04223_),
    .S(1'h1)
  );
  DFFSR _11762_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_0_ ),
    .Q( mem_backbone_0.per_dout_val_0_ ),
    .R(_04224_),
    .S(1'h1)
  );
  DFFSR _11763_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_1_ ),
    .Q( mem_backbone_0.per_dout_val_1_ ),
    .R(_04225_),
    .S(1'h1)
  );
  DFFSR _11764_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_2_ ),
    .Q( mem_backbone_0.per_dout_val_2_ ),
    .R(_04226_),
    .S(1'h1)
  );
  DFFSR _11765_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_3_ ),
    .Q( mem_backbone_0.per_dout_val_3_ ),
    .R(_04227_),
    .S(1'h1)
  );
  DFFSR _11766_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_4_ ),
    .Q( mem_backbone_0.per_dout_val_4_ ),
    .R(_04228_),
    .S(1'h1)
  );
  DFFSR _11767_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_5_ ),
    .Q( mem_backbone_0.per_dout_val_5_ ),
    .R(_04229_),
    .S(1'h1)
  );
  DFFSR _11768_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_6_ ),
    .Q( mem_backbone_0.per_dout_val_6_ ),
    .R(_04230_),
    .S(1'h1)
  );
  DFFSR _11769_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_7_ ),
    .Q( mem_backbone_0.per_dout_val_7_ ),
    .R(_04231_),
    .S(1'h1)
  );
  DFFSR _11770_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_8_ ),
    .Q( mem_backbone_0.per_dout_val_8_ ),
    .R(_04232_),
    .S(1'h1)
  );
  DFFSR _11771_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_9_ ),
    .Q( mem_backbone_0.per_dout_val_9_ ),
    .R(_04233_),
    .S(1'h1)
  );
  DFFSR _11772_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_10_ ),
    .Q( mem_backbone_0.per_dout_val_10_ ),
    .R(_04234_),
    .S(1'h1)
  );
  DFFSR _11773_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_11_ ),
    .Q( mem_backbone_0.per_dout_val_11_ ),
    .R(_04235_),
    .S(1'h1)
  );
  DFFSR _11774_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_12_ ),
    .Q( mem_backbone_0.per_dout_val_12_ ),
    .R(_04236_),
    .S(1'h1)
  );
  DFFSR _11775_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_13_ ),
    .Q( mem_backbone_0.per_dout_val_13_ ),
    .R(_04237_),
    .S(1'h1)
  );
  DFFSR _11776_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_14_ ),
    .Q( mem_backbone_0.per_dout_val_14_ ),
    .R(_04238_),
    .S(1'h1)
  );
  DFFSR _11777_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_15_ ),
    .Q( mem_backbone_0.per_dout_val_15_ ),
    .R(_04239_),
    .S(1'h1)
  );
  INVX1 _11778_ (
    .A( multiplier_0.op1_15_ ),
    .Y(_05298_)
  );
  INVX1 _11779_ (
    .A( multiplier_0.op1_12_ ),
    .Y(_05299_)
  );
  INVX1 _11780_ (
    .A( multiplier_0.op1_8_ ),
    .Y(_05300_)
  );
  INVX1 _11781_ (
    .A( multiplier_0.op1_7_ ),
    .Y(_05301_)
  );
  INVX1 _11782_ (
    .A( multiplier_0.op1_6_ ),
    .Y(_05302_)
  );
  INVX1 _11783_ (
    .A( multiplier_0.op1_5_ ),
    .Y(_05303_)
  );
  INVX1 _11784_ (
    .A( multiplier_0.op1_4_ ),
    .Y(_05304_)
  );
  INVX1 _11785_ (
    .A( multiplier_0.op1_3_ ),
    .Y(_05305_)
  );
  INVX1 _11786_ (
    .A( multiplier_0.op1_2_ ),
    .Y(_05306_)
  );
  INVX1 _11787_ (
    .A( multiplier_0.op1_1_ ),
    .Y(_05307_)
  );
  INVX1 _11788_ (
    .A( multiplier_0.op2_7_ ),
    .Y(_05308_)
  );
  INVX1 _11789_ (
    .A( multiplier_0.op2_6_ ),
    .Y(_05309_)
  );
  INVX1 _11790_ (
    .A( multiplier_0.op2_5_ ),
    .Y(_05310_)
  );
  INVX1 _11791_ (
    .A( multiplier_0.op2_4_ ),
    .Y(_05311_)
  );
  INVX1 _11792_ (
    .A( multiplier_0.op2_3_ ),
    .Y(_05312_)
  );
  INVX1 _11793_ (
    .A( multiplier_0.op2_2_ ),
    .Y(_05313_)
  );
  INVX1 _11794_ (
    .A( multiplier_0.op2_1_ ),
    .Y(_05314_)
  );
  INVX1 _11795_ (
    .A( multiplier_0.op2_0_ ),
    .Y(_05315_)
  );
  INVX1 _11796_ (
    .A( multiplier_0.reslo_15_ ),
    .Y(_05316_)
  );
  INVX1 _11797_ (
    .A( multiplier_0.reslo_13_ ),
    .Y(_05317_)
  );
  INVX1 _11798_ (
    .A( multiplier_0.reslo_10_ ),
    .Y(_05318_)
  );
  INVX1 _11799_ (
    .A( multiplier_0.reslo_2_ ),
    .Y(_05319_)
  );
  INVX1 _11800_ (
    .A( multiplier_0.reslo_0_ ),
    .Y(_05320_)
  );
  INVX1 _11801_ (
    .A( multiplier_0.reshi_13_ ),
    .Y(_05321_)
  );
  INVX1 _11802_ (
    .A( multiplier_0.reshi_12_ ),
    .Y(_05322_)
  );
  INVX1 _11803_ (
    .A( multiplier_0.reshi_11_ ),
    .Y(_05323_)
  );
  INVX1 _11804_ (
    .A( multiplier_0.reshi_9_ ),
    .Y(_05324_)
  );
  INVX1 _11805_ (
    .A( multiplier_0.reshi_8_ ),
    .Y(_05325_)
  );
  INVX1 _11806_ (
    .A( multiplier_0.reshi_5_ ),
    .Y(_05326_)
  );
  INVX1 _11807_ (
    .A( multiplier_0.reshi_4_ ),
    .Y(_05327_)
  );
  INVX1 _11808_ (
    .A( multiplier_0.reshi_3_ ),
    .Y(_05328_)
  );
  INVX1 _11809_ (
    .A( multiplier_0.reshi_2_ ),
    .Y(_05329_)
  );
  INVX1 _11810_ (
    .A( multiplier_0.sumext_10_ ),
    .Y(_05330_)
  );
  INVX1 _11811_ (
    .A( multiplier_0.sumext_0_ ),
    .Y(_05331_)
  );
  INVX1 _11812_ (
    .A( multiplier_0.sign_sel ),
    .Y(_05332_)
  );
  INVX1 _11813_ (
    .A( multiplier_0.cycle_1_ ),
    .Y(_05333_)
  );
  INVX1 _11814_ (
    .A( multiplier_0.cycle_0_ ),
    .Y(_05334_)
  );
  INVX1 _11815_ (
    .A(_06266_),
    .Y(_05335_)
  );
  INVX1 _11816_ (
    .A(_06269_),
    .Y(_05336_)
  );
  INVX1 _11817_ (
    .A(_06271_),
    .Y(_05337_)
  );
  INVX1 _11818_ (
    .A(_06272_),
    .Y(_05338_)
  );
  INVX1 _11819_ (
    .A(_06265_),
    .Y(_05339_)
  );
  INVX1 _11820_ (
    .A(_06327_),
    .Y(_04464_)
  );
  NOR2X1 _11821_ (
    .A(_06293_),
    .B(_06292_),
    .Y(_05340_)
  );
  OR2X1 _11822_ (
    .A(_06264_),
    .B(1'h0),
    .Y(_05341_)
  );
  NAND2X1 _11823_ (
    .A(_05339_),
    .B(_06291_),
    .Y(_05342_)
  );
  NOR2X1 _11824_ (
    .A(_05341_),
    .B(_05342_),
    .Y(_05343_)
  );
  NOR2X1 _11825_ (
    .A(_06273_),
    .B(_05338_),
    .Y(_05344_)
  );
  NOR2X1 _11826_ (
    .A(_06263_),
    .B(_06274_),
    .Y(_05345_)
  );
  NAND2X1 _11827_ (
    .A(_05344_),
    .B(_05345_),
    .Y(_05346_)
  );
  NOR2X1 _11828_ (
    .A(_06271_),
    .B(_06270_),
    .Y(_05347_)
  );
  NAND3X1 _11829_ (
    .A(_06269_),
    .B(_06268_),
    .C(_05347_),
    .Y(_05348_)
  );
  NOR2X1 _11830_ (
    .A(_05346_),
    .B(_05348_),
    .Y(_05349_)
  );
  AND2X1 _11831_ (
    .A(_05343_),
    .B(_05349_),
    .Y(_05350_)
  );
  OAI21X1 _11832_ (
    .A(_06293_),
    .B(_06292_),
    .C(_05350_),
    .Y(_05351_)
  );
  NOR2X1 _11833_ (
    .A(_05338_),
    .B(_06274_),
    .Y(_05352_)
  );
  NAND3X1 _11834_ (
    .A(_06268_),
    .B(_05337_),
    .C(_05352_),
    .Y(_05353_)
  );
  NOR2X1 _11835_ (
    .A(_06273_),
    .B(_06263_),
    .Y(_05354_)
  );
  NOR2X1 _11836_ (
    .A(_05336_),
    .B(_06270_),
    .Y(_05355_)
  );
  NAND3X1 _11837_ (
    .A(_05343_),
    .B(_05354_),
    .C(_05355_),
    .Y(_05356_)
  );
  NOR2X1 _11838_ (
    .A(_05353_),
    .B(_05356_),
    .Y(_05357_)
  );
  OAI21X1 _11839_ (
    .A(_06293_),
    .B(_06292_),
    .C(_05357_),
    .Y(_05358_)
  );
  OR2X1 _11840_ (
    .A(_06267_),
    .B(_05358_),
    .Y(_05359_)
  );
  OAI21X1 _11841_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_15_ ),
    .Y(_05360_)
  );
  AND2X1 _11842_ (
    .A(_06293_),
    .B(_06281_),
    .Y(_05361_)
  );
  NAND2X1 _11843_ (
    .A(_06293_),
    .B(_06281_),
    .Y(_05362_)
  );
  OAI21X1 _11844_ (
    .A(_05359_),
    .B(_05362_),
    .C(_05360_),
    .Y(_04601_)
  );
  OAI21X1 _11845_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_14_ ),
    .Y(_05363_)
  );
  AND2X1 _11846_ (
    .A(_06293_),
    .B(_06280_),
    .Y(_05364_)
  );
  NAND2X1 _11847_ (
    .A(_06293_),
    .B(_06280_),
    .Y(_05365_)
  );
  OAI21X1 _11848_ (
    .A(_05359_),
    .B(_05365_),
    .C(_05363_),
    .Y(_04600_)
  );
  OAI21X1 _11849_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_13_ ),
    .Y(_05366_)
  );
  AND2X1 _11850_ (
    .A(_06293_),
    .B(_06279_),
    .Y(_05367_)
  );
  NAND2X1 _11851_ (
    .A(_06293_),
    .B(_06279_),
    .Y(_05368_)
  );
  OAI21X1 _11852_ (
    .A(_05359_),
    .B(_05368_),
    .C(_05366_),
    .Y(_04599_)
  );
  OAI21X1 _11853_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_12_ ),
    .Y(_05369_)
  );
  AND2X1 _11854_ (
    .A(_06293_),
    .B(_06278_),
    .Y(_05370_)
  );
  NAND2X1 _11855_ (
    .A(_06293_),
    .B(_06278_),
    .Y(_05371_)
  );
  OAI21X1 _11856_ (
    .A(_05359_),
    .B(_05371_),
    .C(_05369_),
    .Y(_04598_)
  );
  OAI21X1 _11857_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_11_ ),
    .Y(_05372_)
  );
  AND2X1 _11858_ (
    .A(_06293_),
    .B(_06277_),
    .Y(_05373_)
  );
  NAND2X1 _11859_ (
    .A(_06293_),
    .B(_06277_),
    .Y(_05374_)
  );
  OAI21X1 _11860_ (
    .A(_05359_),
    .B(_05374_),
    .C(_05372_),
    .Y(_04597_)
  );
  OAI21X1 _11861_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_10_ ),
    .Y(_05375_)
  );
  AND2X1 _11862_ (
    .A(_06293_),
    .B(_06276_),
    .Y(_05376_)
  );
  NAND2X1 _11863_ (
    .A(_06293_),
    .B(_06276_),
    .Y(_05377_)
  );
  OAI21X1 _11864_ (
    .A(_05359_),
    .B(_05377_),
    .C(_05375_),
    .Y(_04596_)
  );
  OAI21X1 _11865_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_9_ ),
    .Y(_05378_)
  );
  AND2X1 _11866_ (
    .A(_06293_),
    .B(_06290_),
    .Y(_05379_)
  );
  NAND2X1 _11867_ (
    .A(_06293_),
    .B(_06290_),
    .Y(_05380_)
  );
  OAI21X1 _11868_ (
    .A(_05359_),
    .B(_05380_),
    .C(_05378_),
    .Y(_04595_)
  );
  OAI21X1 _11869_ (
    .A(_06267_),
    .B(_05351_),
    .C( multiplier_0.op1_8_ ),
    .Y(_05381_)
  );
  AND2X1 _11870_ (
    .A(_06293_),
    .B(_06289_),
    .Y(_05382_)
  );
  NAND2X1 _11871_ (
    .A(_06293_),
    .B(_06289_),
    .Y(_05383_)
  );
  OAI21X1 _11872_ (
    .A(_05359_),
    .B(_05383_),
    .C(_05381_),
    .Y(_04594_)
  );
  MUX2X1 _11873_ (
    .A( multiplier_0.op1_7_ ),
    .B(_06288_),
    .S(_05359_),
    .Y(_05384_)
  );
  INVX1 _11874_ (
    .A(_05384_),
    .Y(_04593_)
  );
  MUX2X1 _11875_ (
    .A( multiplier_0.op1_6_ ),
    .B(_06287_),
    .S(_05359_),
    .Y(_05385_)
  );
  INVX1 _11876_ (
    .A(_05385_),
    .Y(_04592_)
  );
  MUX2X1 _11877_ (
    .A( multiplier_0.op1_5_ ),
    .B(_06286_),
    .S(_05359_),
    .Y(_05386_)
  );
  INVX1 _11878_ (
    .A(_05386_),
    .Y(_04591_)
  );
  MUX2X1 _11879_ (
    .A( multiplier_0.op1_4_ ),
    .B(_06285_),
    .S(_05359_),
    .Y(_05387_)
  );
  INVX1 _11880_ (
    .A(_05387_),
    .Y(_04590_)
  );
  MUX2X1 _11881_ (
    .A( multiplier_0.op1_3_ ),
    .B(_06284_),
    .S(_05359_),
    .Y(_05388_)
  );
  INVX1 _11882_ (
    .A(_05388_),
    .Y(_04589_)
  );
  MUX2X1 _11883_ (
    .A( multiplier_0.op1_2_ ),
    .B(_06283_),
    .S(_05359_),
    .Y(_05389_)
  );
  INVX1 _11884_ (
    .A(_05389_),
    .Y(_04588_)
  );
  MUX2X1 _11885_ (
    .A( multiplier_0.op1_1_ ),
    .B(_06282_),
    .S(_05359_),
    .Y(_05390_)
  );
  INVX1 _11886_ (
    .A(_05390_),
    .Y(_04587_)
  );
  MUX2X1 _11887_ (
    .A( multiplier_0.op1_0_ ),
    .B(_06275_),
    .S(_05359_),
    .Y(_05391_)
  );
  INVX1 _11888_ (
    .A(_05391_),
    .Y(_04586_)
  );
  NAND2X1 _11889_ (
    .A(_06267_),
    .B(_05335_),
    .Y(_05392_)
  );
  OR2X1 _11890_ (
    .A(_06262_),
    .B(_05392_),
    .Y(_05393_)
  );
  NOR2X1 _11891_ (
    .A(_05351_),
    .B(_05393_),
    .Y( multiplier_0.op2_wr )
  );
  OR2X1 _11892_ (
    .A(_05358_),
    .B(_05393_),
    .Y(_05394_)
  );
  OAI21X1 _11893_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_15_ ),
    .Y(_05395_)
  );
  OAI21X1 _11894_ (
    .A(_05362_),
    .B(_05394_),
    .C(_05395_),
    .Y(_04585_)
  );
  OAI21X1 _11895_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_14_ ),
    .Y(_05396_)
  );
  OAI21X1 _11896_ (
    .A(_05365_),
    .B(_05394_),
    .C(_05396_),
    .Y(_04584_)
  );
  OAI21X1 _11897_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_13_ ),
    .Y(_05397_)
  );
  OAI21X1 _11898_ (
    .A(_05368_),
    .B(_05394_),
    .C(_05397_),
    .Y(_04583_)
  );
  OAI21X1 _11899_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_12_ ),
    .Y(_05398_)
  );
  OAI21X1 _11900_ (
    .A(_05371_),
    .B(_05394_),
    .C(_05398_),
    .Y(_04582_)
  );
  OAI21X1 _11901_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_11_ ),
    .Y(_05399_)
  );
  OAI21X1 _11902_ (
    .A(_05374_),
    .B(_05394_),
    .C(_05399_),
    .Y(_04581_)
  );
  OAI21X1 _11903_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_10_ ),
    .Y(_05400_)
  );
  OAI21X1 _11904_ (
    .A(_05377_),
    .B(_05394_),
    .C(_05400_),
    .Y(_04580_)
  );
  OAI21X1 _11905_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_9_ ),
    .Y(_05401_)
  );
  OAI21X1 _11906_ (
    .A(_05380_),
    .B(_05394_),
    .C(_05401_),
    .Y(_04579_)
  );
  OAI21X1 _11907_ (
    .A(_05351_),
    .B(_05393_),
    .C( multiplier_0.op2_8_ ),
    .Y(_05402_)
  );
  OAI21X1 _11908_ (
    .A(_05383_),
    .B(_05394_),
    .C(_05402_),
    .Y(_04578_)
  );
  MUX2X1 _11909_ (
    .A( multiplier_0.op2_7_ ),
    .B(_06288_),
    .S(_05394_),
    .Y(_05403_)
  );
  INVX1 _11910_ (
    .A(_05403_),
    .Y(_04577_)
  );
  MUX2X1 _11911_ (
    .A( multiplier_0.op2_6_ ),
    .B(_06287_),
    .S(_05394_),
    .Y(_05404_)
  );
  INVX1 _11912_ (
    .A(_05404_),
    .Y(_04576_)
  );
  MUX2X1 _11913_ (
    .A( multiplier_0.op2_5_ ),
    .B(_06286_),
    .S(_05394_),
    .Y(_05405_)
  );
  INVX1 _11914_ (
    .A(_05405_),
    .Y(_04575_)
  );
  MUX2X1 _11915_ (
    .A( multiplier_0.op2_4_ ),
    .B(_06285_),
    .S(_05394_),
    .Y(_05406_)
  );
  INVX1 _11916_ (
    .A(_05406_),
    .Y(_04574_)
  );
  MUX2X1 _11917_ (
    .A( multiplier_0.op2_3_ ),
    .B(_06284_),
    .S(_05394_),
    .Y(_05407_)
  );
  INVX1 _11918_ (
    .A(_05407_),
    .Y(_04573_)
  );
  MUX2X1 _11919_ (
    .A( multiplier_0.op2_2_ ),
    .B(_06283_),
    .S(_05394_),
    .Y(_05408_)
  );
  INVX1 _11920_ (
    .A(_05408_),
    .Y(_04572_)
  );
  MUX2X1 _11921_ (
    .A( multiplier_0.op2_1_ ),
    .B(_06282_),
    .S(_05394_),
    .Y(_05409_)
  );
  INVX1 _11922_ (
    .A(_05409_),
    .Y(_04571_)
  );
  MUX2X1 _11923_ (
    .A( multiplier_0.op2_0_ ),
    .B(_06275_),
    .S(_05394_),
    .Y(_05410_)
  );
  INVX1 _11924_ (
    .A(_05410_),
    .Y(_04570_)
  );
  NOR2X1 _11925_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05411_)
  );
  NAND2X1 _11926_ (
    .A(_05333_),
    .B(_05334_),
    .Y(_05412_)
  );
  NAND3X1 _11927_ (
    .A(_06267_),
    .B(_05335_),
    .C(_06262_),
    .Y(_05413_)
  );
  NOR2X1 _11928_ (
    .A(_05351_),
    .B(_05413_),
    .Y(_05414_)
  );
  OAI22X1 _11929_ (
    .A( multiplier_0.acc_sel ),
    .B(_05394_),
    .C(_05413_),
    .D(_05358_),
    .Y(_05415_)
  );
  NOR2X1 _11930_ (
    .A(_05412_),
    .B(_05415_),
    .Y(_05416_)
  );
  OR2X1 _11931_ (
    .A(_05412_),
    .B(_05415_),
    .Y(_05417_)
  );
  NAND2X1 _11932_ (
    .A( multiplier_0.op2_9_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05418_)
  );
  MUX2X1 _11933_ (
    .A( multiplier_0.op2_9_ ),
    .B( multiplier_0.op2_1_ ),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05419_)
  );
  OAI21X1 _11934_ (
    .A(_05314_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05418_),
    .Y(_05420_)
  );
  NAND2X1 _11935_ (
    .A( multiplier_0.op2_8_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05421_)
  );
  MUX2X1 _11936_ (
    .A( multiplier_0.op2_8_ ),
    .B( multiplier_0.op2_0_ ),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05422_)
  );
  OAI21X1 _11937_ (
    .A(_05315_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05421_),
    .Y(_05423_)
  );
  NAND2X1 _11938_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05423_),
    .Y(_05424_)
  );
  NAND2X1 _11939_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05420_),
    .Y(_05425_)
  );
  OR2X1 _11940_ (
    .A(_05300_),
    .B(_05422_),
    .Y(_05426_)
  );
  NOR2X1 _11941_ (
    .A(_05425_),
    .B(_05426_),
    .Y(_05427_)
  );
  NAND2X1 _11942_ (
    .A( multiplier_0.op2_10_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05428_)
  );
  OAI21X1 _11943_ (
    .A(_05313_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05428_),
    .Y(_05429_)
  );
  NAND2X1 _11944_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05429_),
    .Y(_05430_)
  );
  OAI21X1 _11945_ (
    .A(_05300_),
    .B(_05419_),
    .C(_05424_),
    .Y(_05431_)
  );
  OAI21X1 _11946_ (
    .A(_05425_),
    .B(_05426_),
    .C(_05431_),
    .Y(_05432_)
  );
  NOR2X1 _11947_ (
    .A(_05430_),
    .B(_05432_),
    .Y(_05433_)
  );
  NOR2X1 _11948_ (
    .A(_05427_),
    .B(_05433_),
    .Y(_05434_)
  );
  NAND2X1 _11949_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05429_),
    .Y(_05435_)
  );
  NAND2X1 _11950_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05423_),
    .Y(_05436_)
  );
  AND2X1 _11951_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05420_),
    .Y(_05437_)
  );
  XNOR2X1 _11952_ (
    .A(_05425_),
    .B(_05436_),
    .Y(_05438_)
  );
  NAND2X1 _11953_ (
    .A(_05435_),
    .B(_05438_),
    .Y(_05439_)
  );
  OR2X1 _11954_ (
    .A(_05435_),
    .B(_05438_),
    .Y(_05440_)
  );
  NAND2X1 _11955_ (
    .A(_05439_),
    .B(_05440_),
    .Y(_05441_)
  );
  NOR2X1 _11956_ (
    .A(_05434_),
    .B(_05441_),
    .Y(_05442_)
  );
  NAND2X1 _11957_ (
    .A( multiplier_0.op2_13_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05443_)
  );
  OAI21X1 _11958_ (
    .A(_05310_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05443_),
    .Y(_05444_)
  );
  NAND2X1 _11959_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05444_),
    .Y(_05445_)
  );
  NAND2X1 _11960_ (
    .A( multiplier_0.op2_12_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05446_)
  );
  OAI21X1 _11961_ (
    .A(_05311_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05446_),
    .Y(_05447_)
  );
  NAND2X1 _11962_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05447_),
    .Y(_05448_)
  );
  NAND2X1 _11963_ (
    .A( multiplier_0.op2_11_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05449_)
  );
  OAI21X1 _11964_ (
    .A(_05312_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05449_),
    .Y(_05450_)
  );
  NAND2X1 _11965_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05450_),
    .Y(_05451_)
  );
  NAND2X1 _11966_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05447_),
    .Y(_05452_)
  );
  NAND2X1 _11967_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05450_),
    .Y(_05453_)
  );
  XNOR2X1 _11968_ (
    .A(_05448_),
    .B(_05451_),
    .Y(_05454_)
  );
  XNOR2X1 _11969_ (
    .A(_05445_),
    .B(_05454_),
    .Y(_05455_)
  );
  INVX1 _11970_ (
    .A(_05455_),
    .Y(_05456_)
  );
  XOR2X1 _11971_ (
    .A(_05434_),
    .B(_05441_),
    .Y(_05457_)
  );
  AOI21X1 _11972_ (
    .A(_05456_),
    .B(_05457_),
    .C(_05442_),
    .Y(_05458_)
  );
  INVX1 _11973_ (
    .A(_05458_),
    .Y(_05459_)
  );
  NAND2X1 _11974_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05444_),
    .Y(_05460_)
  );
  NAND2X1 _11975_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05450_),
    .Y(_05461_)
  );
  AND2X1 _11976_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05447_),
    .Y(_05462_)
  );
  OR2X1 _11977_ (
    .A(_05452_),
    .B(_05461_),
    .Y(_05463_)
  );
  XNOR2X1 _11978_ (
    .A(_05452_),
    .B(_05461_),
    .Y(_05464_)
  );
  XNOR2X1 _11979_ (
    .A(_05460_),
    .B(_05464_),
    .Y(_05465_)
  );
  OAI21X1 _11980_ (
    .A(_05425_),
    .B(_05436_),
    .C(_05440_),
    .Y(_05466_)
  );
  NAND2X1 _11981_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05429_),
    .Y(_05467_)
  );
  NAND2X1 _11982_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05423_),
    .Y(_05468_)
  );
  AND2X1 _11983_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05420_),
    .Y(_05469_)
  );
  NAND3X1 _11984_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05423_),
    .C(_05437_),
    .Y(_05470_)
  );
  XOR2X1 _11985_ (
    .A(_05437_),
    .B(_05468_),
    .Y(_05471_)
  );
  XNOR2X1 _11986_ (
    .A(_05467_),
    .B(_05471_),
    .Y(_05472_)
  );
  INVX1 _11987_ (
    .A(_05472_),
    .Y(_05473_)
  );
  NAND2X1 _11988_ (
    .A(_05466_),
    .B(_05473_),
    .Y(_05474_)
  );
  XNOR2X1 _11989_ (
    .A(_05466_),
    .B(_05473_),
    .Y(_05475_)
  );
  XOR2X1 _11990_ (
    .A(_05465_),
    .B(_05475_),
    .Y(_05476_)
  );
  NAND2X1 _11991_ (
    .A(_05459_),
    .B(_05476_),
    .Y(_05477_)
  );
  NAND2X1 _11992_ (
    .A( multiplier_0.op2_15_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05478_)
  );
  OAI21X1 _11993_ (
    .A(_05308_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05478_),
    .Y(_05479_)
  );
  NAND2X1 _11994_ (
    .A( multiplier_0.op2_14_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_05480_)
  );
  OAI21X1 _11995_ (
    .A(_05309_),
    .B( multiplier_0.cycle_0_ ),
    .C(_05480_),
    .Y(_05481_)
  );
  INVX1 _11996_ (
    .A(_05481_),
    .Y(_05482_)
  );
  NAND2X1 _11997_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05479_),
    .Y(_05483_)
  );
  NAND2X1 _11998_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05481_),
    .Y(_05484_)
  );
  OR2X1 _11999_ (
    .A(_05332_),
    .B(_05478_),
    .Y(_05485_)
  );
  NOR2X1 _12000_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05485_),
    .Y(_05486_)
  );
  INVX1 _12001_ (
    .A(_05486_),
    .Y(_05487_)
  );
  AOI22X1 _12002_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05479_),
    .C(_05481_),
    .D( multiplier_0.op1_4_ ),
    .Y(_05488_)
  );
  INVX1 _12003_ (
    .A(_05488_),
    .Y(_05489_)
  );
  OAI21X1 _12004_ (
    .A(_05483_),
    .B(_05484_),
    .C(_05489_),
    .Y(_05490_)
  );
  OAI22X1 _12005_ (
    .A(_05483_),
    .B(_05484_),
    .C(_05487_),
    .D(_05490_),
    .Y(_05491_)
  );
  NOR2X1 _12006_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05485_),
    .Y(_05492_)
  );
  INVX1 _12007_ (
    .A(_05492_),
    .Y(_05493_)
  );
  AND2X1 _12008_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05479_),
    .Y(_05494_)
  );
  NAND3X1 _12009_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05481_),
    .C(_05494_),
    .Y(_05495_)
  );
  OAI21X1 _12010_ (
    .A(_05303_),
    .B(_05482_),
    .C(_05483_),
    .Y(_05496_)
  );
  NAND2X1 _12011_ (
    .A(_05495_),
    .B(_05496_),
    .Y(_05497_)
  );
  XNOR2X1 _12012_ (
    .A(_05493_),
    .B(_05497_),
    .Y(_05498_)
  );
  INVX1 _12013_ (
    .A(_05498_),
    .Y(_05499_)
  );
  OAI22X1 _12014_ (
    .A(_05452_),
    .B(_05453_),
    .C(_05454_),
    .D(_05445_),
    .Y(_05500_)
  );
  NAND2X1 _12015_ (
    .A(_05499_),
    .B(_05500_),
    .Y(_05501_)
  );
  XOR2X1 _12016_ (
    .A(_05498_),
    .B(_05500_),
    .Y(_05502_)
  );
  INVX1 _12017_ (
    .A(_05502_),
    .Y(_05503_)
  );
  NAND2X1 _12018_ (
    .A(_05491_),
    .B(_05503_),
    .Y(_05504_)
  );
  XOR2X1 _12019_ (
    .A(_05491_),
    .B(_05502_),
    .Y(_05505_)
  );
  NOR2X1 _12020_ (
    .A(_05459_),
    .B(_05476_),
    .Y(_05506_)
  );
  XNOR2X1 _12021_ (
    .A(_05458_),
    .B(_05476_),
    .Y(_05507_)
  );
  OAI21X1 _12022_ (
    .A(_05505_),
    .B(_05506_),
    .C(_05477_),
    .Y(_05508_)
  );
  OAI21X1 _12023_ (
    .A(_05493_),
    .B(_05497_),
    .C(_05495_),
    .Y(_05509_)
  );
  NOR2X1 _12024_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05485_),
    .Y(_05510_)
  );
  INVX1 _12025_ (
    .A(_05510_),
    .Y(_05511_)
  );
  NAND2X1 _12026_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05481_),
    .Y(_05512_)
  );
  NAND2X1 _12027_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05479_),
    .Y(_05513_)
  );
  NAND3X1 _12028_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05481_),
    .C(_05494_),
    .Y(_05514_)
  );
  XOR2X1 _12029_ (
    .A(_05494_),
    .B(_05512_),
    .Y(_05515_)
  );
  XNOR2X1 _12030_ (
    .A(_05511_),
    .B(_05515_),
    .Y(_05516_)
  );
  OAI21X1 _12031_ (
    .A(_05460_),
    .B(_05464_),
    .C(_05463_),
    .Y(_05517_)
  );
  INVX1 _12032_ (
    .A(_05517_),
    .Y(_05518_)
  );
  XOR2X1 _12033_ (
    .A(_05516_),
    .B(_05517_),
    .Y(_05519_)
  );
  INVX1 _12034_ (
    .A(_05519_),
    .Y(_05520_)
  );
  NAND2X1 _12035_ (
    .A(_05509_),
    .B(_05520_),
    .Y(_05521_)
  );
  XOR2X1 _12036_ (
    .A(_05509_),
    .B(_05519_),
    .Y(_05522_)
  );
  OAI21X1 _12037_ (
    .A(_05465_),
    .B(_05475_),
    .C(_05474_),
    .Y(_05523_)
  );
  NAND2X1 _12038_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05444_),
    .Y(_05524_)
  );
  NAND2X1 _12039_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05450_),
    .Y(_05525_)
  );
  AND2X1 _12040_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05447_),
    .Y(_05526_)
  );
  NAND3X1 _12041_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05450_),
    .C(_05462_),
    .Y(_05527_)
  );
  XOR2X1 _12042_ (
    .A(_05462_),
    .B(_05525_),
    .Y(_05528_)
  );
  XNOR2X1 _12043_ (
    .A(_05524_),
    .B(_05528_),
    .Y(_05529_)
  );
  OAI21X1 _12044_ (
    .A(_05467_),
    .B(_05471_),
    .C(_05470_),
    .Y(_05530_)
  );
  NAND2X1 _12045_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05429_),
    .Y(_05531_)
  );
  NAND2X1 _12046_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05423_),
    .Y(_05532_)
  );
  NAND3X1 _12047_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05423_),
    .C(_05469_),
    .Y(_05533_)
  );
  XOR2X1 _12048_ (
    .A(_05469_),
    .B(_05532_),
    .Y(_05534_)
  );
  XNOR2X1 _12049_ (
    .A(_05531_),
    .B(_05534_),
    .Y(_05535_)
  );
  INVX1 _12050_ (
    .A(_05535_),
    .Y(_05536_)
  );
  NAND2X1 _12051_ (
    .A(_05530_),
    .B(_05536_),
    .Y(_05537_)
  );
  XOR2X1 _12052_ (
    .A(_05530_),
    .B(_05535_),
    .Y(_05538_)
  );
  XOR2X1 _12053_ (
    .A(_05529_),
    .B(_05538_),
    .Y(_05539_)
  );
  NAND2X1 _12054_ (
    .A(_05523_),
    .B(_05539_),
    .Y(_05540_)
  );
  XNOR2X1 _12055_ (
    .A(_05523_),
    .B(_05539_),
    .Y(_05541_)
  );
  XOR2X1 _12056_ (
    .A(_05522_),
    .B(_05541_),
    .Y(_05542_)
  );
  NAND2X1 _12057_ (
    .A(_05508_),
    .B(_05542_),
    .Y(_05543_)
  );
  AND2X1 _12058_ (
    .A(_05501_),
    .B(_05504_),
    .Y(_05544_)
  );
  XNOR2X1 _12059_ (
    .A(_05508_),
    .B(_05542_),
    .Y(_05545_)
  );
  OAI21X1 _12060_ (
    .A(_05544_),
    .B(_05545_),
    .C(_05543_),
    .Y(_05546_)
  );
  OAI21X1 _12061_ (
    .A(_05516_),
    .B(_05518_),
    .C(_05521_),
    .Y(_05547_)
  );
  INVX1 _12062_ (
    .A(_05547_),
    .Y(_05548_)
  );
  OAI21X1 _12063_ (
    .A(_05522_),
    .B(_05541_),
    .C(_05540_),
    .Y(_05549_)
  );
  OAI21X1 _12064_ (
    .A(_05511_),
    .B(_05515_),
    .C(_05514_),
    .Y(_05550_)
  );
  NOR2X1 _12065_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05485_),
    .Y(_05551_)
  );
  INVX1 _12066_ (
    .A(_05551_),
    .Y(_05552_)
  );
  NAND2X1 _12067_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05481_),
    .Y(_05553_)
  );
  NAND2X1 _12068_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05479_),
    .Y(_05554_)
  );
  OAI21X1 _12069_ (
    .A(_05301_),
    .B(_05482_),
    .C(_05513_),
    .Y(_05555_)
  );
  OAI21X1 _12070_ (
    .A(_05512_),
    .B(_05554_),
    .C(_05555_),
    .Y(_05556_)
  );
  XNOR2X1 _12071_ (
    .A(_05552_),
    .B(_05556_),
    .Y(_05557_)
  );
  OAI21X1 _12072_ (
    .A(_05524_),
    .B(_05528_),
    .C(_05527_),
    .Y(_05558_)
  );
  INVX1 _12073_ (
    .A(_05558_),
    .Y(_05559_)
  );
  XOR2X1 _12074_ (
    .A(_05557_),
    .B(_05558_),
    .Y(_05560_)
  );
  INVX1 _12075_ (
    .A(_05560_),
    .Y(_05561_)
  );
  NAND2X1 _12076_ (
    .A(_05550_),
    .B(_05561_),
    .Y(_05562_)
  );
  XOR2X1 _12077_ (
    .A(_05550_),
    .B(_05560_),
    .Y(_05563_)
  );
  OAI21X1 _12078_ (
    .A(_05529_),
    .B(_05538_),
    .C(_05537_),
    .Y(_05564_)
  );
  NAND2X1 _12079_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05444_),
    .Y(_05565_)
  );
  NAND2X1 _12080_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05450_),
    .Y(_05566_)
  );
  AND2X1 _12081_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05447_),
    .Y(_05567_)
  );
  NAND3X1 _12082_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05450_),
    .C(_05526_),
    .Y(_05568_)
  );
  XOR2X1 _12083_ (
    .A(_05526_),
    .B(_05566_),
    .Y(_05569_)
  );
  XNOR2X1 _12084_ (
    .A(_05565_),
    .B(_05569_),
    .Y(_05570_)
  );
  OAI21X1 _12085_ (
    .A(_05531_),
    .B(_05534_),
    .C(_05533_),
    .Y(_05571_)
  );
  NAND2X1 _12086_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05429_),
    .Y(_05572_)
  );
  NAND2X1 _12087_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05423_),
    .Y(_05573_)
  );
  NAND2X1 _12088_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05420_),
    .Y(_05574_)
  );
  OAI21X1 _12089_ (
    .A(_05299_),
    .B(_05419_),
    .C(_05573_),
    .Y(_05575_)
  );
  OAI21X1 _12090_ (
    .A(_05532_),
    .B(_05574_),
    .C(_05575_),
    .Y(_05576_)
  );
  XNOR2X1 _12091_ (
    .A(_05572_),
    .B(_05576_),
    .Y(_05577_)
  );
  INVX1 _12092_ (
    .A(_05577_),
    .Y(_05578_)
  );
  NAND2X1 _12093_ (
    .A(_05571_),
    .B(_05578_),
    .Y(_05579_)
  );
  XOR2X1 _12094_ (
    .A(_05571_),
    .B(_05577_),
    .Y(_05580_)
  );
  XOR2X1 _12095_ (
    .A(_05570_),
    .B(_05580_),
    .Y(_05581_)
  );
  NAND2X1 _12096_ (
    .A(_05564_),
    .B(_05581_),
    .Y(_05582_)
  );
  XNOR2X1 _12097_ (
    .A(_05564_),
    .B(_05581_),
    .Y(_05583_)
  );
  XOR2X1 _12098_ (
    .A(_05563_),
    .B(_05583_),
    .Y(_05584_)
  );
  NAND2X1 _12099_ (
    .A(_05549_),
    .B(_05584_),
    .Y(_05585_)
  );
  XNOR2X1 _12100_ (
    .A(_05549_),
    .B(_05584_),
    .Y(_05586_)
  );
  XNOR2X1 _12101_ (
    .A(_05547_),
    .B(_05586_),
    .Y(_05587_)
  );
  NAND2X1 _12102_ (
    .A(_05546_),
    .B(_05587_),
    .Y(_05588_)
  );
  OAI21X1 _12103_ (
    .A(_05548_),
    .B(_05586_),
    .C(_05585_),
    .Y(_05589_)
  );
  OAI21X1 _12104_ (
    .A(_05557_),
    .B(_05559_),
    .C(_05562_),
    .Y(_05590_)
  );
  INVX1 _12105_ (
    .A(_05590_),
    .Y(_05591_)
  );
  OAI21X1 _12106_ (
    .A(_05563_),
    .B(_05583_),
    .C(_05582_),
    .Y(_05592_)
  );
  OAI22X1 _12107_ (
    .A(_05512_),
    .B(_05554_),
    .C(_05556_),
    .D(_05552_),
    .Y(_05593_)
  );
  NOR2X1 _12108_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05485_),
    .Y(_05594_)
  );
  INVX1 _12109_ (
    .A(_05594_),
    .Y(_05595_)
  );
  NAND2X1 _12110_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05481_),
    .Y(_05596_)
  );
  NAND2X1 _12111_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05479_),
    .Y(_05597_)
  );
  OAI21X1 _12112_ (
    .A(_05300_),
    .B(_05482_),
    .C(_05554_),
    .Y(_05598_)
  );
  OAI21X1 _12113_ (
    .A(_05553_),
    .B(_05597_),
    .C(_05598_),
    .Y(_05599_)
  );
  XNOR2X1 _12114_ (
    .A(_05595_),
    .B(_05599_),
    .Y(_05600_)
  );
  OAI21X1 _12115_ (
    .A(_05565_),
    .B(_05569_),
    .C(_05568_),
    .Y(_05601_)
  );
  INVX1 _12116_ (
    .A(_05601_),
    .Y(_05602_)
  );
  XOR2X1 _12117_ (
    .A(_05600_),
    .B(_05601_),
    .Y(_05603_)
  );
  INVX1 _12118_ (
    .A(_05603_),
    .Y(_05604_)
  );
  NAND2X1 _12119_ (
    .A(_05593_),
    .B(_05604_),
    .Y(_05605_)
  );
  XOR2X1 _12120_ (
    .A(_05593_),
    .B(_05603_),
    .Y(_05606_)
  );
  OAI21X1 _12121_ (
    .A(_05570_),
    .B(_05580_),
    .C(_05579_),
    .Y(_05607_)
  );
  NAND2X1 _12122_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05444_),
    .Y(_05608_)
  );
  NAND2X1 _12123_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05450_),
    .Y(_05609_)
  );
  AND2X1 _12124_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05447_),
    .Y(_05610_)
  );
  NAND3X1 _12125_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05450_),
    .C(_05567_),
    .Y(_05611_)
  );
  XOR2X1 _12126_ (
    .A(_05567_),
    .B(_05609_),
    .Y(_05612_)
  );
  XNOR2X1 _12127_ (
    .A(_05608_),
    .B(_05612_),
    .Y(_05613_)
  );
  OAI22X1 _12128_ (
    .A(_05532_),
    .B(_05574_),
    .C(_05576_),
    .D(_05572_),
    .Y(_05614_)
  );
  NAND2X1 _12129_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05429_),
    .Y(_05615_)
  );
  NAND2X1 _12130_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05423_),
    .Y(_05616_)
  );
  NAND2X1 _12131_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05420_),
    .Y(_05617_)
  );
  NAND2X1 _12132_ (
    .A(_05574_),
    .B(_05616_),
    .Y(_05618_)
  );
  OAI21X1 _12133_ (
    .A(_05573_),
    .B(_05617_),
    .C(_05618_),
    .Y(_05619_)
  );
  XNOR2X1 _12134_ (
    .A(_05615_),
    .B(_05619_),
    .Y(_05620_)
  );
  INVX1 _12135_ (
    .A(_05620_),
    .Y(_05621_)
  );
  NAND2X1 _12136_ (
    .A(_05614_),
    .B(_05621_),
    .Y(_05622_)
  );
  XOR2X1 _12137_ (
    .A(_05614_),
    .B(_05620_),
    .Y(_05623_)
  );
  XOR2X1 _12138_ (
    .A(_05613_),
    .B(_05623_),
    .Y(_05624_)
  );
  NAND2X1 _12139_ (
    .A(_05607_),
    .B(_05624_),
    .Y(_05625_)
  );
  XNOR2X1 _12140_ (
    .A(_05607_),
    .B(_05624_),
    .Y(_05626_)
  );
  XOR2X1 _12141_ (
    .A(_05606_),
    .B(_05626_),
    .Y(_05627_)
  );
  NAND2X1 _12142_ (
    .A(_05592_),
    .B(_05627_),
    .Y(_05628_)
  );
  XNOR2X1 _12143_ (
    .A(_05592_),
    .B(_05627_),
    .Y(_05629_)
  );
  XNOR2X1 _12144_ (
    .A(_05590_),
    .B(_05629_),
    .Y(_05630_)
  );
  NAND2X1 _12145_ (
    .A(_05589_),
    .B(_05630_),
    .Y(_05631_)
  );
  XNOR2X1 _12146_ (
    .A(_05589_),
    .B(_05630_),
    .Y(_05632_)
  );
  NOR2X1 _12147_ (
    .A(_05588_),
    .B(_05632_),
    .Y(_05633_)
  );
  XOR2X1 _12148_ (
    .A(_05588_),
    .B(_05632_),
    .Y(_05634_)
  );
  NOR2X1 _12149_ (
    .A(_05426_),
    .B(_05485_),
    .Y(_05635_)
  );
  OR2X1 _12150_ (
    .A(_05301_),
    .B(_05419_),
    .Y(_05636_)
  );
  XNOR2X1 _12151_ (
    .A(_05426_),
    .B(_05485_),
    .Y(_05637_)
  );
  NOR2X1 _12152_ (
    .A(_05636_),
    .B(_05637_),
    .Y(_05638_)
  );
  NOR2X1 _12153_ (
    .A(_05635_),
    .B(_05638_),
    .Y(_05639_)
  );
  XNOR2X1 _12154_ (
    .A(_05430_),
    .B(_05432_),
    .Y(_05640_)
  );
  OR2X1 _12155_ (
    .A(_05639_),
    .B(_05640_),
    .Y(_05641_)
  );
  NAND2X1 _12156_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05444_),
    .Y(_05642_)
  );
  NAND2X1 _12157_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05447_),
    .Y(_05643_)
  );
  NAND2X1 _12158_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05450_),
    .Y(_05644_)
  );
  XNOR2X1 _12159_ (
    .A(_05453_),
    .B(_05643_),
    .Y(_05645_)
  );
  XNOR2X1 _12160_ (
    .A(_05642_),
    .B(_05645_),
    .Y(_05646_)
  );
  XNOR2X1 _12161_ (
    .A(_05639_),
    .B(_05640_),
    .Y(_05647_)
  );
  OAI21X1 _12162_ (
    .A(_05646_),
    .B(_05647_),
    .C(_05641_),
    .Y(_05648_)
  );
  XNOR2X1 _12163_ (
    .A(_05455_),
    .B(_05457_),
    .Y(_05649_)
  );
  NAND2X1 _12164_ (
    .A(_05648_),
    .B(_05649_),
    .Y(_05650_)
  );
  NAND2X1 _12165_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05479_),
    .Y(_05651_)
  );
  NAND2X1 _12166_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05481_),
    .Y(_05652_)
  );
  OR2X1 _12167_ (
    .A(_05484_),
    .B(_05651_),
    .Y(_05653_)
  );
  NOR2X1 _12168_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05485_),
    .Y(_05654_)
  );
  OAI21X1 _12169_ (
    .A(_05305_),
    .B(_05482_),
    .C(_05651_),
    .Y(_05655_)
  );
  NAND2X1 _12170_ (
    .A(_05653_),
    .B(_05655_),
    .Y(_05656_)
  );
  NAND3X1 _12171_ (
    .A(_05653_),
    .B(_05654_),
    .C(_05655_),
    .Y(_05657_)
  );
  OAI21X1 _12172_ (
    .A(_05484_),
    .B(_05651_),
    .C(_05657_),
    .Y(_05658_)
  );
  XNOR2X1 _12173_ (
    .A(_05487_),
    .B(_05490_),
    .Y(_05659_)
  );
  INVX1 _12174_ (
    .A(_05659_),
    .Y(_05660_)
  );
  OAI22X1 _12175_ (
    .A(_05448_),
    .B(_05644_),
    .C(_05645_),
    .D(_05642_),
    .Y(_05661_)
  );
  XOR2X1 _12176_ (
    .A(_05659_),
    .B(_05661_),
    .Y(_05662_)
  );
  AOI21X1 _12177_ (
    .A(_05653_),
    .B(_05657_),
    .C(_05662_),
    .Y(_05663_)
  );
  XOR2X1 _12178_ (
    .A(_05658_),
    .B(_05662_),
    .Y(_05664_)
  );
  XNOR2X1 _12179_ (
    .A(_05648_),
    .B(_05649_),
    .Y(_05665_)
  );
  OAI21X1 _12180_ (
    .A(_05664_),
    .B(_05665_),
    .C(_05650_),
    .Y(_05666_)
  );
  XNOR2X1 _12181_ (
    .A(_05505_),
    .B(_05507_),
    .Y(_05667_)
  );
  NAND2X1 _12182_ (
    .A(_05666_),
    .B(_05667_),
    .Y(_05668_)
  );
  AOI21X1 _12183_ (
    .A(_05660_),
    .B(_05661_),
    .C(_05663_),
    .Y(_05669_)
  );
  XNOR2X1 _12184_ (
    .A(_05666_),
    .B(_05667_),
    .Y(_05670_)
  );
  OAI21X1 _12185_ (
    .A(_05669_),
    .B(_05670_),
    .C(_05668_),
    .Y(_05671_)
  );
  XOR2X1 _12186_ (
    .A(_05544_),
    .B(_05545_),
    .Y(_05672_)
  );
  NAND2X1 _12187_ (
    .A(_05671_),
    .B(_05672_),
    .Y(_05673_)
  );
  XNOR2X1 _12188_ (
    .A(_05546_),
    .B(_05587_),
    .Y(_05674_)
  );
  AND2X1 _12189_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05675_)
  );
  NOR2X1 _12190_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05676_)
  );
  OR2X1 _12191_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05677_)
  );
  NOR2X1 _12192_ (
    .A(_05302_),
    .B(_05422_),
    .Y(_05678_)
  );
  OR2X1 _12193_ (
    .A(_05302_),
    .B(_05422_),
    .Y(_05679_)
  );
  NOR2X1 _12194_ (
    .A(_05636_),
    .B(_05679_),
    .Y(_05680_)
  );
  AND2X1 _12195_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05429_),
    .Y(_05681_)
  );
  OAI22X1 _12196_ (
    .A(_05302_),
    .B(_05419_),
    .C(_05422_),
    .D(_05301_),
    .Y(_05682_)
  );
  OAI21X1 _12197_ (
    .A(_05636_),
    .B(_05679_),
    .C(_05682_),
    .Y(_05683_)
  );
  AOI21X1 _12198_ (
    .A(_05681_),
    .B(_05682_),
    .C(_05680_),
    .Y(_05684_)
  );
  XNOR2X1 _12199_ (
    .A(_05636_),
    .B(_05637_),
    .Y(_05685_)
  );
  NAND2X1 _12200_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05447_),
    .Y(_05686_)
  );
  NAND2X1 _12201_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05429_),
    .Y(_05687_)
  );
  XNOR2X1 _12202_ (
    .A(_05644_),
    .B(_05687_),
    .Y(_05688_)
  );
  OR2X1 _12203_ (
    .A(_05686_),
    .B(_05688_),
    .Y(_05689_)
  );
  XNOR2X1 _12204_ (
    .A(_05686_),
    .B(_05688_),
    .Y(_05690_)
  );
  INVX1 _12205_ (
    .A(_05690_),
    .Y(_05691_)
  );
  XOR2X1 _12206_ (
    .A(_05684_),
    .B(_05685_),
    .Y(_05692_)
  );
  NAND2X1 _12207_ (
    .A(_05691_),
    .B(_05692_),
    .Y(_05693_)
  );
  OAI21X1 _12208_ (
    .A(_05684_),
    .B(_05685_),
    .C(_05693_),
    .Y(_05694_)
  );
  XOR2X1 _12209_ (
    .A(_05646_),
    .B(_05647_),
    .Y(_05695_)
  );
  NAND2X1 _12210_ (
    .A(_05694_),
    .B(_05695_),
    .Y(_05696_)
  );
  NAND2X1 _12211_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05444_),
    .Y(_05697_)
  );
  NAND2X1 _12212_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05444_),
    .Y(_05698_)
  );
  NAND2X1 _12213_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05479_),
    .Y(_05699_)
  );
  XNOR2X1 _12214_ (
    .A(_05652_),
    .B(_05697_),
    .Y(_05700_)
  );
  OAI22X1 _12215_ (
    .A(_05484_),
    .B(_05698_),
    .C(_05699_),
    .D(_05700_),
    .Y(_05701_)
  );
  XOR2X1 _12216_ (
    .A(_05654_),
    .B(_05656_),
    .Y(_05702_)
  );
  INVX1 _12217_ (
    .A(_05702_),
    .Y(_05703_)
  );
  OAI21X1 _12218_ (
    .A(_05644_),
    .B(_05687_),
    .C(_05689_),
    .Y(_05704_)
  );
  NAND2X1 _12219_ (
    .A(_05703_),
    .B(_05704_),
    .Y(_05705_)
  );
  XOR2X1 _12220_ (
    .A(_05702_),
    .B(_05704_),
    .Y(_05706_)
  );
  INVX1 _12221_ (
    .A(_05706_),
    .Y(_05707_)
  );
  NAND2X1 _12222_ (
    .A(_05701_),
    .B(_05707_),
    .Y(_05708_)
  );
  XOR2X1 _12223_ (
    .A(_05701_),
    .B(_05706_),
    .Y(_05709_)
  );
  XNOR2X1 _12224_ (
    .A(_05694_),
    .B(_05695_),
    .Y(_05710_)
  );
  OAI21X1 _12225_ (
    .A(_05709_),
    .B(_05710_),
    .C(_05696_),
    .Y(_05711_)
  );
  XOR2X1 _12226_ (
    .A(_05664_),
    .B(_05665_),
    .Y(_05712_)
  );
  NAND2X1 _12227_ (
    .A(_05711_),
    .B(_05712_),
    .Y(_05713_)
  );
  AND2X1 _12228_ (
    .A(_05705_),
    .B(_05708_),
    .Y(_05714_)
  );
  XNOR2X1 _12229_ (
    .A(_05711_),
    .B(_05712_),
    .Y(_05715_)
  );
  OAI21X1 _12230_ (
    .A(_05714_),
    .B(_05715_),
    .C(_05713_),
    .Y(_05716_)
  );
  XOR2X1 _12231_ (
    .A(_05669_),
    .B(_05670_),
    .Y(_05717_)
  );
  NAND2X1 _12232_ (
    .A(_05716_),
    .B(_05717_),
    .Y(_05718_)
  );
  XNOR2X1 _12233_ (
    .A(_05671_),
    .B(_05672_),
    .Y(_05719_)
  );
  NOR2X1 _12234_ (
    .A(_05718_),
    .B(_05719_),
    .Y(_05720_)
  );
  XOR2X1 _12235_ (
    .A(_05718_),
    .B(_05719_),
    .Y(_05721_)
  );
  NOR2X1 _12236_ (
    .A(_05303_),
    .B(_05419_),
    .Y(_05722_)
  );
  NOR2X1 _12237_ (
    .A(_05303_),
    .B(_05422_),
    .Y(_05723_)
  );
  NAND2X1 _12238_ (
    .A(_05678_),
    .B(_05722_),
    .Y(_05724_)
  );
  NAND2X1 _12239_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05429_),
    .Y(_05725_)
  );
  NOR2X1 _12240_ (
    .A(_05678_),
    .B(_05722_),
    .Y(_05726_)
  );
  XNOR2X1 _12241_ (
    .A(_05679_),
    .B(_05722_),
    .Y(_05727_)
  );
  OAI21X1 _12242_ (
    .A(_05725_),
    .B(_05726_),
    .C(_05724_),
    .Y(_05728_)
  );
  XNOR2X1 _12243_ (
    .A(_05681_),
    .B(_05683_),
    .Y(_05729_)
  );
  NAND2X1 _12244_ (
    .A(_05728_),
    .B(_05729_),
    .Y(_05730_)
  );
  NAND2X1 _12245_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05447_),
    .Y(_05731_)
  );
  NAND2X1 _12246_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05450_),
    .Y(_05732_)
  );
  NAND2X1 _12247_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05450_),
    .Y(_05733_)
  );
  XNOR2X1 _12248_ (
    .A(_05731_),
    .B(_05732_),
    .Y(_05734_)
  );
  XNOR2X1 _12249_ (
    .A(_05698_),
    .B(_05734_),
    .Y(_05735_)
  );
  XNOR2X1 _12250_ (
    .A(_05728_),
    .B(_05729_),
    .Y(_05736_)
  );
  OAI21X1 _12251_ (
    .A(_05735_),
    .B(_05736_),
    .C(_05730_),
    .Y(_05737_)
  );
  XNOR2X1 _12252_ (
    .A(_05690_),
    .B(_05692_),
    .Y(_05738_)
  );
  NAND2X1 _12253_ (
    .A(_05737_),
    .B(_05738_),
    .Y(_05739_)
  );
  AND2X1 _12254_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05481_),
    .Y(_05740_)
  );
  NAND3X1 _12255_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05479_),
    .C(_05740_),
    .Y(_05741_)
  );
  INVX1 _12256_ (
    .A(_05741_),
    .Y(_05742_)
  );
  XNOR2X1 _12257_ (
    .A(_05699_),
    .B(_05700_),
    .Y(_05743_)
  );
  INVX1 _12258_ (
    .A(_05743_),
    .Y(_05744_)
  );
  OAI22X1 _12259_ (
    .A(_05686_),
    .B(_05733_),
    .C(_05734_),
    .D(_05698_),
    .Y(_05745_)
  );
  XOR2X1 _12260_ (
    .A(_05743_),
    .B(_05745_),
    .Y(_05746_)
  );
  NOR2X1 _12261_ (
    .A(_05741_),
    .B(_05746_),
    .Y(_05747_)
  );
  XNOR2X1 _12262_ (
    .A(_05741_),
    .B(_05746_),
    .Y(_05748_)
  );
  XNOR2X1 _12263_ (
    .A(_05737_),
    .B(_05738_),
    .Y(_05749_)
  );
  OAI21X1 _12264_ (
    .A(_05748_),
    .B(_05749_),
    .C(_05739_),
    .Y(_05750_)
  );
  XOR2X1 _12265_ (
    .A(_05709_),
    .B(_05710_),
    .Y(_05751_)
  );
  NAND2X1 _12266_ (
    .A(_05750_),
    .B(_05751_),
    .Y(_05752_)
  );
  AOI21X1 _12267_ (
    .A(_05744_),
    .B(_05745_),
    .C(_05747_),
    .Y(_05753_)
  );
  XNOR2X1 _12268_ (
    .A(_05750_),
    .B(_05751_),
    .Y(_05754_)
  );
  OAI21X1 _12269_ (
    .A(_05753_),
    .B(_05754_),
    .C(_05752_),
    .Y(_05755_)
  );
  XOR2X1 _12270_ (
    .A(_05714_),
    .B(_05715_),
    .Y(_05756_)
  );
  NAND2X1 _12271_ (
    .A(_05755_),
    .B(_05756_),
    .Y(_05757_)
  );
  XNOR2X1 _12272_ (
    .A(_05716_),
    .B(_05717_),
    .Y(_05758_)
  );
  OR2X1 _12273_ (
    .A(_05757_),
    .B(_05758_),
    .Y(_05759_)
  );
  XOR2X1 _12274_ (
    .A(_05757_),
    .B(_05758_),
    .Y(_05760_)
  );
  INVX1 _12275_ (
    .A(_05760_),
    .Y(_05761_)
  );
  NOR2X1 _12276_ (
    .A(_05304_),
    .B(_05419_),
    .Y(_05762_)
  );
  NOR2X1 _12277_ (
    .A(_05304_),
    .B(_05422_),
    .Y(_05763_)
  );
  NAND2X1 _12278_ (
    .A(_05723_),
    .B(_05762_),
    .Y(_05764_)
  );
  NAND2X1 _12279_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05429_),
    .Y(_05765_)
  );
  XNOR2X1 _12280_ (
    .A(_05723_),
    .B(_05762_),
    .Y(_05766_)
  );
  OAI21X1 _12281_ (
    .A(_05765_),
    .B(_05766_),
    .C(_05764_),
    .Y(_05767_)
  );
  XNOR2X1 _12282_ (
    .A(_05725_),
    .B(_05727_),
    .Y(_05768_)
  );
  NAND2X1 _12283_ (
    .A(_05767_),
    .B(_05768_),
    .Y(_05769_)
  );
  NAND2X1 _12284_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05444_),
    .Y(_05770_)
  );
  NAND2X1 _12285_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05447_),
    .Y(_05771_)
  );
  AND2X1 _12286_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05450_),
    .Y(_05772_)
  );
  OR2X1 _12287_ (
    .A(_05733_),
    .B(_05771_),
    .Y(_05773_)
  );
  XNOR2X1 _12288_ (
    .A(_05733_),
    .B(_05771_),
    .Y(_05774_)
  );
  XNOR2X1 _12289_ (
    .A(_05770_),
    .B(_05774_),
    .Y(_05775_)
  );
  XNOR2X1 _12290_ (
    .A(_05767_),
    .B(_05768_),
    .Y(_05776_)
  );
  OAI21X1 _12291_ (
    .A(_05775_),
    .B(_05776_),
    .C(_05769_),
    .Y(_05777_)
  );
  XOR2X1 _12292_ (
    .A(_05735_),
    .B(_05736_),
    .Y(_05778_)
  );
  NAND2X1 _12293_ (
    .A(_05777_),
    .B(_05778_),
    .Y(_05779_)
  );
  AOI22X1 _12294_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05479_),
    .C(_05481_),
    .D( multiplier_0.op1_1_ ),
    .Y(_05780_)
  );
  NOR2X1 _12295_ (
    .A(_05742_),
    .B(_05780_),
    .Y(_05781_)
  );
  OAI21X1 _12296_ (
    .A(_05770_),
    .B(_05774_),
    .C(_05773_),
    .Y(_05782_)
  );
  NAND2X1 _12297_ (
    .A(_05781_),
    .B(_05782_),
    .Y(_05783_)
  );
  XNOR2X1 _12298_ (
    .A(_05781_),
    .B(_05782_),
    .Y(_05784_)
  );
  XNOR2X1 _12299_ (
    .A(_05777_),
    .B(_05778_),
    .Y(_05785_)
  );
  OAI21X1 _12300_ (
    .A(_05784_),
    .B(_05785_),
    .C(_05779_),
    .Y(_05786_)
  );
  XNOR2X1 _12301_ (
    .A(_05748_),
    .B(_05749_),
    .Y(_05787_)
  );
  INVX1 _12302_ (
    .A(_05787_),
    .Y(_05788_)
  );
  NAND2X1 _12303_ (
    .A(_05786_),
    .B(_05788_),
    .Y(_05789_)
  );
  XOR2X1 _12304_ (
    .A(_05786_),
    .B(_05787_),
    .Y(_05790_)
  );
  OAI21X1 _12305_ (
    .A(_05783_),
    .B(_05790_),
    .C(_05789_),
    .Y(_05791_)
  );
  XNOR2X1 _12306_ (
    .A(_05753_),
    .B(_05754_),
    .Y(_05792_)
  );
  INVX1 _12307_ (
    .A(_05792_),
    .Y(_05793_)
  );
  NAND2X1 _12308_ (
    .A(_05791_),
    .B(_05793_),
    .Y(_05794_)
  );
  XNOR2X1 _12309_ (
    .A(_05755_),
    .B(_05756_),
    .Y(_05795_)
  );
  NOR2X1 _12310_ (
    .A(_05794_),
    .B(_05795_),
    .Y(_05796_)
  );
  XOR2X1 _12311_ (
    .A(_05794_),
    .B(_05795_),
    .Y(_05797_)
  );
  NOR2X1 _12312_ (
    .A(_05305_),
    .B(_05419_),
    .Y(_05798_)
  );
  NOR2X1 _12313_ (
    .A(_05305_),
    .B(_05422_),
    .Y(_05799_)
  );
  NAND2X1 _12314_ (
    .A(_05763_),
    .B(_05798_),
    .Y(_05800_)
  );
  NAND2X1 _12315_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05429_),
    .Y(_05801_)
  );
  XNOR2X1 _12316_ (
    .A(_05763_),
    .B(_05798_),
    .Y(_05802_)
  );
  OAI21X1 _12317_ (
    .A(_05801_),
    .B(_05802_),
    .C(_05800_),
    .Y(_05803_)
  );
  XOR2X1 _12318_ (
    .A(_05765_),
    .B(_05766_),
    .Y(_05804_)
  );
  NAND2X1 _12319_ (
    .A(_05803_),
    .B(_05804_),
    .Y(_05805_)
  );
  NAND2X1 _12320_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05444_),
    .Y(_05806_)
  );
  NAND2X1 _12321_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05447_),
    .Y(_05807_)
  );
  NAND3X1 _12322_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05447_),
    .C(_05772_),
    .Y(_05808_)
  );
  XOR2X1 _12323_ (
    .A(_05772_),
    .B(_05807_),
    .Y(_05809_)
  );
  XNOR2X1 _12324_ (
    .A(_05806_),
    .B(_05809_),
    .Y(_05810_)
  );
  XNOR2X1 _12325_ (
    .A(_05803_),
    .B(_05804_),
    .Y(_05811_)
  );
  OAI21X1 _12326_ (
    .A(_05810_),
    .B(_05811_),
    .C(_05805_),
    .Y(_05812_)
  );
  XOR2X1 _12327_ (
    .A(_05775_),
    .B(_05776_),
    .Y(_05813_)
  );
  NAND2X1 _12328_ (
    .A(_05812_),
    .B(_05813_),
    .Y(_05814_)
  );
  OAI21X1 _12329_ (
    .A(_05806_),
    .B(_05809_),
    .C(_05808_),
    .Y(_05815_)
  );
  NAND2X1 _12330_ (
    .A(_05740_),
    .B(_05815_),
    .Y(_05816_)
  );
  XNOR2X1 _12331_ (
    .A(_05740_),
    .B(_05815_),
    .Y(_05817_)
  );
  XNOR2X1 _12332_ (
    .A(_05812_),
    .B(_05813_),
    .Y(_05818_)
  );
  OAI21X1 _12333_ (
    .A(_05817_),
    .B(_05818_),
    .C(_05814_),
    .Y(_05819_)
  );
  XOR2X1 _12334_ (
    .A(_05784_),
    .B(_05785_),
    .Y(_05820_)
  );
  NAND2X1 _12335_ (
    .A(_05819_),
    .B(_05820_),
    .Y(_05821_)
  );
  XNOR2X1 _12336_ (
    .A(_05819_),
    .B(_05820_),
    .Y(_05822_)
  );
  OAI21X1 _12337_ (
    .A(_05816_),
    .B(_05822_),
    .C(_05821_),
    .Y(_05823_)
  );
  XOR2X1 _12338_ (
    .A(_05783_),
    .B(_05790_),
    .Y(_05824_)
  );
  OR2X1 _12339_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05485_),
    .Y(_05825_)
  );
  XNOR2X1 _12340_ (
    .A(_05823_),
    .B(_05824_),
    .Y(_05826_)
  );
  NOR2X1 _12341_ (
    .A(_05825_),
    .B(_05826_),
    .Y(_05827_)
  );
  AOI21X1 _12342_ (
    .A(_05823_),
    .B(_05824_),
    .C(_05827_),
    .Y(_05828_)
  );
  XOR2X1 _12343_ (
    .A(_05791_),
    .B(_05792_),
    .Y(_05829_)
  );
  OR2X1 _12344_ (
    .A(_05828_),
    .B(_05829_),
    .Y(_05830_)
  );
  XNOR2X1 _12345_ (
    .A(_05828_),
    .B(_05829_),
    .Y(_05831_)
  );
  OR2X1 _12346_ (
    .A(_05306_),
    .B(_05419_),
    .Y(_05832_)
  );
  NAND3X1 _12347_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05420_),
    .C(_05799_),
    .Y(_05833_)
  );
  NAND2X1 _12348_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05429_),
    .Y(_05834_)
  );
  XOR2X1 _12349_ (
    .A(_05799_),
    .B(_05832_),
    .Y(_05835_)
  );
  OAI21X1 _12350_ (
    .A(_05834_),
    .B(_05835_),
    .C(_05833_),
    .Y(_05836_)
  );
  XOR2X1 _12351_ (
    .A(_05801_),
    .B(_05802_),
    .Y(_05837_)
  );
  NAND2X1 _12352_ (
    .A(_05836_),
    .B(_05837_),
    .Y(_05838_)
  );
  NAND2X1 _12353_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05450_),
    .Y(_05839_)
  );
  NOR2X1 _12354_ (
    .A(_05807_),
    .B(_05839_),
    .Y(_05840_)
  );
  OR2X1 _12355_ (
    .A(_05807_),
    .B(_05839_),
    .Y(_05841_)
  );
  AOI22X1 _12356_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05447_),
    .C(_05450_),
    .D( multiplier_0.op1_1_ ),
    .Y(_05842_)
  );
  OR2X1 _12357_ (
    .A(_05840_),
    .B(_05842_),
    .Y(_05843_)
  );
  XNOR2X1 _12358_ (
    .A(_05836_),
    .B(_05837_),
    .Y(_05844_)
  );
  OAI21X1 _12359_ (
    .A(_05843_),
    .B(_05844_),
    .C(_05838_),
    .Y(_05845_)
  );
  XOR2X1 _12360_ (
    .A(_05810_),
    .B(_05811_),
    .Y(_05846_)
  );
  NAND2X1 _12361_ (
    .A(_05845_),
    .B(_05846_),
    .Y(_05847_)
  );
  XNOR2X1 _12362_ (
    .A(_05845_),
    .B(_05846_),
    .Y(_05848_)
  );
  OAI21X1 _12363_ (
    .A(_05841_),
    .B(_05848_),
    .C(_05847_),
    .Y(_05849_)
  );
  XOR2X1 _12364_ (
    .A(_05817_),
    .B(_05818_),
    .Y(_05850_)
  );
  NAND2X1 _12365_ (
    .A(_05849_),
    .B(_05850_),
    .Y(_05851_)
  );
  XNOR2X1 _12366_ (
    .A(_05816_),
    .B(_05822_),
    .Y(_05852_)
  );
  OR2X1 _12367_ (
    .A(_05851_),
    .B(_05852_),
    .Y(_05853_)
  );
  XNOR2X1 _12368_ (
    .A(_05825_),
    .B(_05826_),
    .Y(_05854_)
  );
  NOR2X1 _12369_ (
    .A(_05853_),
    .B(_05854_),
    .Y(_05855_)
  );
  NOR2X1 _12370_ (
    .A(_05307_),
    .B(_05422_),
    .Y(_05856_)
  );
  OR2X1 _12371_ (
    .A(_05307_),
    .B(_05422_),
    .Y(_05857_)
  );
  NAND2X1 _12372_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05429_),
    .Y(_05858_)
  );
  OAI22X1 _12373_ (
    .A(_05307_),
    .B(_05419_),
    .C(_05422_),
    .D(_05306_),
    .Y(_05859_)
  );
  OAI21X1 _12374_ (
    .A(_05832_),
    .B(_05857_),
    .C(_05859_),
    .Y(_05860_)
  );
  OAI22X1 _12375_ (
    .A(_05832_),
    .B(_05857_),
    .C(_05858_),
    .D(_05860_),
    .Y(_05861_)
  );
  XOR2X1 _12376_ (
    .A(_05834_),
    .B(_05835_),
    .Y(_05862_)
  );
  NAND2X1 _12377_ (
    .A(_05861_),
    .B(_05862_),
    .Y(_05863_)
  );
  XNOR2X1 _12378_ (
    .A(_05861_),
    .B(_05862_),
    .Y(_05864_)
  );
  OAI21X1 _12379_ (
    .A(_05839_),
    .B(_05864_),
    .C(_05863_),
    .Y(_05865_)
  );
  XOR2X1 _12380_ (
    .A(_05843_),
    .B(_05844_),
    .Y(_05866_)
  );
  NAND2X1 _12381_ (
    .A(_05865_),
    .B(_05866_),
    .Y(_05867_)
  );
  XNOR2X1 _12382_ (
    .A(_05841_),
    .B(_05848_),
    .Y(_05868_)
  );
  OR2X1 _12383_ (
    .A(_05867_),
    .B(_05868_),
    .Y(_05869_)
  );
  XNOR2X1 _12384_ (
    .A(_05849_),
    .B(_05850_),
    .Y(_05870_)
  );
  NOR2X1 _12385_ (
    .A(_05869_),
    .B(_05870_),
    .Y(_05871_)
  );
  XOR2X1 _12386_ (
    .A(_05851_),
    .B(_05852_),
    .Y(_05872_)
  );
  NAND2X1 _12387_ (
    .A(_05871_),
    .B(_05872_),
    .Y(_05873_)
  );
  NAND3X1 _12388_ (
    .A( multiplier_0.op1_0_ ),
    .B( multiplier_0.op2_0_ ),
    .C(_05334_),
    .Y(_05874_)
  );
  NAND2X1 _12389_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05420_),
    .Y(_05875_)
  );
  OR2X1 _12390_ (
    .A(_05857_),
    .B(_05875_),
    .Y(_05876_)
  );
  XNOR2X1 _12391_ (
    .A(_05858_),
    .B(_05860_),
    .Y(_05877_)
  );
  NOR2X1 _12392_ (
    .A(_05876_),
    .B(_05877_),
    .Y(_05878_)
  );
  INVX1 _12393_ (
    .A(_05878_),
    .Y(_05879_)
  );
  XNOR2X1 _12394_ (
    .A(_05839_),
    .B(_05864_),
    .Y(_05880_)
  );
  OR2X1 _12395_ (
    .A(_05879_),
    .B(_05880_),
    .Y(_05881_)
  );
  XNOR2X1 _12396_ (
    .A(_05865_),
    .B(_05866_),
    .Y(_05882_)
  );
  NOR2X1 _12397_ (
    .A(_05881_),
    .B(_05882_),
    .Y(_05883_)
  );
  XOR2X1 _12398_ (
    .A(_05867_),
    .B(_05868_),
    .Y(_05884_)
  );
  NAND2X1 _12399_ (
    .A(_05883_),
    .B(_05884_),
    .Y(_05885_)
  );
  XNOR2X1 _12400_ (
    .A(_05869_),
    .B(_05870_),
    .Y(_05886_)
  );
  NOR2X1 _12401_ (
    .A(_05885_),
    .B(_05886_),
    .Y(_05887_)
  );
  INVX1 _12402_ (
    .A(_05887_),
    .Y(_05888_)
  );
  XNOR2X1 _12403_ (
    .A(_05871_),
    .B(_05872_),
    .Y(_05889_)
  );
  OAI21X1 _12404_ (
    .A(_05888_),
    .B(_05889_),
    .C(_05873_),
    .Y(_05890_)
  );
  XOR2X1 _12405_ (
    .A(_05853_),
    .B(_05854_),
    .Y(_05891_)
  );
  AOI21X1 _12406_ (
    .A(_05890_),
    .B(_05891_),
    .C(_05855_),
    .Y(_05892_)
  );
  OAI21X1 _12407_ (
    .A(_05831_),
    .B(_05892_),
    .C(_05830_),
    .Y(_05893_)
  );
  AOI21X1 _12408_ (
    .A(_05797_),
    .B(_05893_),
    .C(_05796_),
    .Y(_05894_)
  );
  OAI21X1 _12409_ (
    .A(_05761_),
    .B(_05894_),
    .C(_05759_),
    .Y(_05895_)
  );
  AOI21X1 _12410_ (
    .A(_05721_),
    .B(_05895_),
    .C(_05720_),
    .Y(_05896_)
  );
  NOR2X1 _12411_ (
    .A(_05675_),
    .B(_05676_),
    .Y(_05897_)
  );
  OAI21X1 _12412_ (
    .A(_05675_),
    .B(_05896_),
    .C(_05677_),
    .Y(_05898_)
  );
  XNOR2X1 _12413_ (
    .A(_05634_),
    .B(_05898_),
    .Y(_05899_)
  );
  XOR2X1 _12414_ (
    .A(_05885_),
    .B(_05886_),
    .Y(_05900_)
  );
  NAND2X1 _12415_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05900_),
    .Y(_05901_)
  );
  OAI21X1 _12416_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05899_),
    .C(_05901_),
    .Y(_05902_)
  );
  NAND2X1 _12417_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_05902_),
    .Y(_05903_)
  );
  XNOR2X1 _12418_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_05902_),
    .Y(_05904_)
  );
  XNOR2X1 _12419_ (
    .A(_05896_),
    .B(_05897_),
    .Y(_05905_)
  );
  XNOR2X1 _12420_ (
    .A(_05883_),
    .B(_05884_),
    .Y(_05906_)
  );
  NAND2X1 _12421_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05906_),
    .Y(_05907_)
  );
  OAI21X1 _12422_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05905_),
    .C(_05907_),
    .Y(_05908_)
  );
  NOR2X1 _12423_ (
    .A(_05317_),
    .B(_05908_),
    .Y(_05909_)
  );
  XNOR2X1 _12424_ (
    .A( multiplier_0.reslo_13_ ),
    .B(_05908_),
    .Y(_05910_)
  );
  XNOR2X1 _12425_ (
    .A(_05721_),
    .B(_05895_),
    .Y(_05911_)
  );
  XNOR2X1 _12426_ (
    .A(_05881_),
    .B(_05882_),
    .Y(_05912_)
  );
  MUX2X1 _12427_ (
    .A(_05911_),
    .B(_05912_),
    .S(_05334_),
    .Y(_05913_)
  );
  NAND2X1 _12428_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_05913_),
    .Y(_05914_)
  );
  XNOR2X1 _12429_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_05913_),
    .Y(_05915_)
  );
  XNOR2X1 _12430_ (
    .A(_05761_),
    .B(_05894_),
    .Y(_05916_)
  );
  XNOR2X1 _12431_ (
    .A(_05878_),
    .B(_05880_),
    .Y(_05917_)
  );
  NAND2X1 _12432_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05917_),
    .Y(_05918_)
  );
  OAI21X1 _12433_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05916_),
    .C(_05918_),
    .Y(_05919_)
  );
  AND2X1 _12434_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_05919_),
    .Y(_05920_)
  );
  NAND2X1 _12435_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_05919_),
    .Y(_05921_)
  );
  OR2X1 _12436_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_05919_),
    .Y(_05922_)
  );
  NAND2X1 _12437_ (
    .A(_05921_),
    .B(_05922_),
    .Y(_05923_)
  );
  XOR2X1 _12438_ (
    .A(_05797_),
    .B(_05893_),
    .Y(_05924_)
  );
  OAI21X1 _12439_ (
    .A(_05857_),
    .B(_05875_),
    .C(_05877_),
    .Y(_05925_)
  );
  NAND2X1 _12440_ (
    .A(_05879_),
    .B(_05925_),
    .Y(_05926_)
  );
  NAND2X1 _12441_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05926_),
    .Y(_05927_)
  );
  OAI21X1 _12442_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05924_),
    .C(_05927_),
    .Y(_05928_)
  );
  OR2X1 _12443_ (
    .A(_05318_),
    .B(_05928_),
    .Y(_05929_)
  );
  XNOR2X1 _12444_ (
    .A(_05318_),
    .B(_05928_),
    .Y(_05930_)
  );
  XNOR2X1 _12445_ (
    .A(_05831_),
    .B(_05892_),
    .Y(_05931_)
  );
  XNOR2X1 _12446_ (
    .A(_05856_),
    .B(_05875_),
    .Y(_05932_)
  );
  NAND2X1 _12447_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05932_),
    .Y(_05933_)
  );
  OAI21X1 _12448_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05931_),
    .C(_05933_),
    .Y(_05934_)
  );
  AND2X1 _12449_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_05934_),
    .Y(_05935_)
  );
  NAND2X1 _12450_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_05934_),
    .Y(_05936_)
  );
  OR2X1 _12451_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_05934_),
    .Y(_05937_)
  );
  NAND2X1 _12452_ (
    .A(_05936_),
    .B(_05937_),
    .Y(_05938_)
  );
  XNOR2X1 _12453_ (
    .A(_05890_),
    .B(_05891_),
    .Y(_05939_)
  );
  AOI21X1 _12454_ (
    .A( multiplier_0.op1_0_ ),
    .B( multiplier_0.op2_8_ ),
    .C(_05334_),
    .Y(_05940_)
  );
  AOI21X1 _12455_ (
    .A(_05334_),
    .B(_05939_),
    .C(_05940_),
    .Y(_05941_)
  );
  NAND2X1 _12456_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_05941_),
    .Y(_05942_)
  );
  XNOR2X1 _12457_ (
    .A(_05888_),
    .B(_05889_),
    .Y(_05943_)
  );
  NOR2X1 _12458_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05943_),
    .Y(_05944_)
  );
  AND2X1 _12459_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_05944_),
    .Y(_05945_)
  );
  NAND2X1 _12460_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_05944_),
    .Y(_05946_)
  );
  OR2X1 _12461_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_05944_),
    .Y(_05947_)
  );
  NAND2X1 _12462_ (
    .A(_05946_),
    .B(_05947_),
    .Y(_05948_)
  );
  NAND2X1 _12463_ (
    .A(_05334_),
    .B(_05900_),
    .Y(_05949_)
  );
  NAND3X1 _12464_ (
    .A( multiplier_0.reslo_6_ ),
    .B(_05334_),
    .C(_05900_),
    .Y(_05950_)
  );
  AOI21X1 _12465_ (
    .A(_05334_),
    .B(_05900_),
    .C( multiplier_0.reslo_6_ ),
    .Y(_05951_)
  );
  XNOR2X1 _12466_ (
    .A( multiplier_0.reslo_6_ ),
    .B(_05949_),
    .Y(_05952_)
  );
  NOR2X1 _12467_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05906_),
    .Y(_05953_)
  );
  NAND2X1 _12468_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_05953_),
    .Y(_05954_)
  );
  INVX1 _12469_ (
    .A(_05954_),
    .Y(_05955_)
  );
  OR2X1 _12470_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_05953_),
    .Y(_05956_)
  );
  NAND2X1 _12471_ (
    .A(_05954_),
    .B(_05956_),
    .Y(_05957_)
  );
  NOR2X1 _12472_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05912_),
    .Y(_05958_)
  );
  NAND2X1 _12473_ (
    .A( multiplier_0.reslo_4_ ),
    .B(_05958_),
    .Y(_05959_)
  );
  NAND2X1 _12474_ (
    .A(_05334_),
    .B(_05917_),
    .Y(_05960_)
  );
  NAND3X1 _12475_ (
    .A( multiplier_0.reslo_3_ ),
    .B(_05334_),
    .C(_05917_),
    .Y(_05961_)
  );
  AOI21X1 _12476_ (
    .A(_05334_),
    .B(_05917_),
    .C( multiplier_0.reslo_3_ ),
    .Y(_05962_)
  );
  XNOR2X1 _12477_ (
    .A( multiplier_0.reslo_3_ ),
    .B(_05960_),
    .Y(_05963_)
  );
  NOR2X1 _12478_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05926_),
    .Y(_05964_)
  );
  AND2X1 _12479_ (
    .A( multiplier_0.reslo_2_ ),
    .B(_05964_),
    .Y(_05965_)
  );
  XNOR2X1 _12480_ (
    .A(_05319_),
    .B(_05964_),
    .Y(_05966_)
  );
  AND2X1 _12481_ (
    .A(_05334_),
    .B(_05932_),
    .Y(_05967_)
  );
  NAND2X1 _12482_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_05967_),
    .Y(_05968_)
  );
  NOR2X1 _12483_ (
    .A(_05320_),
    .B(_05874_),
    .Y(_05969_)
  );
  INVX1 _12484_ (
    .A(_05969_),
    .Y(_05970_)
  );
  NOR2X1 _12485_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_05967_),
    .Y(_05971_)
  );
  XOR2X1 _12486_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_05967_),
    .Y(_05972_)
  );
  OAI21X1 _12487_ (
    .A(_05970_),
    .B(_05971_),
    .C(_05968_),
    .Y(_05973_)
  );
  AOI21X1 _12488_ (
    .A(_05966_),
    .B(_05973_),
    .C(_05965_),
    .Y(_05974_)
  );
  OAI21X1 _12489_ (
    .A(_05962_),
    .B(_05974_),
    .C(_05961_),
    .Y(_05975_)
  );
  XOR2X1 _12490_ (
    .A( multiplier_0.reslo_4_ ),
    .B(_05958_),
    .Y(_05976_)
  );
  NAND2X1 _12491_ (
    .A(_05975_),
    .B(_05976_),
    .Y(_05977_)
  );
  NAND2X1 _12492_ (
    .A(_05959_),
    .B(_05977_),
    .Y(_05978_)
  );
  AOI21X1 _12493_ (
    .A(_05956_),
    .B(_05978_),
    .C(_05955_),
    .Y(_05979_)
  );
  OAI21X1 _12494_ (
    .A(_05951_),
    .B(_05979_),
    .C(_05950_),
    .Y(_05980_)
  );
  AOI21X1 _12495_ (
    .A(_05947_),
    .B(_05980_),
    .C(_05945_),
    .Y(_05981_)
  );
  XNOR2X1 _12496_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_05941_),
    .Y(_05982_)
  );
  OAI21X1 _12497_ (
    .A(_05981_),
    .B(_05982_),
    .C(_05942_),
    .Y(_05983_)
  );
  AOI21X1 _12498_ (
    .A(_05937_),
    .B(_05983_),
    .C(_05935_),
    .Y(_05984_)
  );
  OAI21X1 _12499_ (
    .A(_05930_),
    .B(_05984_),
    .C(_05929_),
    .Y(_05985_)
  );
  AOI21X1 _12500_ (
    .A(_05922_),
    .B(_05985_),
    .C(_05920_),
    .Y(_05986_)
  );
  OAI21X1 _12501_ (
    .A(_05915_),
    .B(_05986_),
    .C(_05914_),
    .Y(_05987_)
  );
  AOI21X1 _12502_ (
    .A(_05910_),
    .B(_05987_),
    .C(_05909_),
    .Y(_05988_)
  );
  OR2X1 _12503_ (
    .A(_05904_),
    .B(_05988_),
    .Y(_05989_)
  );
  OAI21X1 _12504_ (
    .A(_05904_),
    .B(_05988_),
    .C(_05903_),
    .Y(_05990_)
  );
  OAI21X1 _12505_ (
    .A(_05591_),
    .B(_05629_),
    .C(_05628_),
    .Y(_05991_)
  );
  OAI21X1 _12506_ (
    .A(_05600_),
    .B(_05602_),
    .C(_05605_),
    .Y(_05992_)
  );
  INVX1 _12507_ (
    .A(_05992_),
    .Y(_05993_)
  );
  OAI21X1 _12508_ (
    .A(_05606_),
    .B(_05626_),
    .C(_05625_),
    .Y(_05994_)
  );
  OAI22X1 _12509_ (
    .A(_05553_),
    .B(_05597_),
    .C(_05599_),
    .D(_05595_),
    .Y(_05995_)
  );
  NOR2X1 _12510_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05485_),
    .Y(_05996_)
  );
  INVX1 _12511_ (
    .A(_05996_),
    .Y(_05997_)
  );
  NAND2X1 _12512_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05481_),
    .Y(_05998_)
  );
  NAND2X1 _12513_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05479_),
    .Y(_05999_)
  );
  NAND2X1 _12514_ (
    .A(_05597_),
    .B(_05998_),
    .Y(_06000_)
  );
  OAI21X1 _12515_ (
    .A(_05596_),
    .B(_05999_),
    .C(_06000_),
    .Y(_06001_)
  );
  XNOR2X1 _12516_ (
    .A(_05997_),
    .B(_06001_),
    .Y(_06002_)
  );
  OAI21X1 _12517_ (
    .A(_05608_),
    .B(_05612_),
    .C(_05611_),
    .Y(_06003_)
  );
  INVX1 _12518_ (
    .A(_06003_),
    .Y(_04602_)
  );
  XOR2X1 _12519_ (
    .A(_06002_),
    .B(_06003_),
    .Y(_04603_)
  );
  INVX1 _12520_ (
    .A(_04603_),
    .Y(_04604_)
  );
  NAND2X1 _12521_ (
    .A(_05995_),
    .B(_04604_),
    .Y(_04605_)
  );
  XOR2X1 _12522_ (
    .A(_05995_),
    .B(_04603_),
    .Y(_04606_)
  );
  OAI21X1 _12523_ (
    .A(_05613_),
    .B(_05623_),
    .C(_05622_),
    .Y(_04607_)
  );
  NAND2X1 _12524_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05444_),
    .Y(_04608_)
  );
  NAND2X1 _12525_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05450_),
    .Y(_04609_)
  );
  NAND2X1 _12526_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05447_),
    .Y(_04610_)
  );
  OR2X1 _12527_ (
    .A(_05609_),
    .B(_04610_),
    .Y(_04611_)
  );
  XOR2X1 _12528_ (
    .A(_05610_),
    .B(_04609_),
    .Y(_04612_)
  );
  XNOR2X1 _12529_ (
    .A(_04608_),
    .B(_04612_),
    .Y(_04613_)
  );
  OAI22X1 _12530_ (
    .A(_05573_),
    .B(_05617_),
    .C(_05619_),
    .D(_05615_),
    .Y(_04614_)
  );
  NAND2X1 _12531_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05429_),
    .Y(_04615_)
  );
  NAND2X1 _12532_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05420_),
    .Y(_04616_)
  );
  INVX1 _12533_ (
    .A(_04616_),
    .Y(_04617_)
  );
  OAI21X1 _12534_ (
    .A(_05298_),
    .B(_05422_),
    .C(_05617_),
    .Y(_04618_)
  );
  OAI21X1 _12535_ (
    .A(_05616_),
    .B(_04616_),
    .C(_04618_),
    .Y(_04619_)
  );
  XNOR2X1 _12536_ (
    .A(_04615_),
    .B(_04619_),
    .Y(_04620_)
  );
  INVX1 _12537_ (
    .A(_04620_),
    .Y(_04621_)
  );
  NAND2X1 _12538_ (
    .A(_04614_),
    .B(_04621_),
    .Y(_04622_)
  );
  XOR2X1 _12539_ (
    .A(_04614_),
    .B(_04620_),
    .Y(_04623_)
  );
  XOR2X1 _12540_ (
    .A(_04613_),
    .B(_04623_),
    .Y(_04624_)
  );
  NAND2X1 _12541_ (
    .A(_04607_),
    .B(_04624_),
    .Y(_04625_)
  );
  XNOR2X1 _12542_ (
    .A(_04607_),
    .B(_04624_),
    .Y(_04626_)
  );
  XOR2X1 _12543_ (
    .A(_04606_),
    .B(_04626_),
    .Y(_04627_)
  );
  NAND2X1 _12544_ (
    .A(_05994_),
    .B(_04627_),
    .Y(_04628_)
  );
  XNOR2X1 _12545_ (
    .A(_05994_),
    .B(_04627_),
    .Y(_04629_)
  );
  XNOR2X1 _12546_ (
    .A(_05992_),
    .B(_04629_),
    .Y(_04630_)
  );
  NAND2X1 _12547_ (
    .A(_05991_),
    .B(_04630_),
    .Y(_04631_)
  );
  XNOR2X1 _12548_ (
    .A(_05991_),
    .B(_04630_),
    .Y(_04632_)
  );
  OR2X1 _12549_ (
    .A(_05631_),
    .B(_04632_),
    .Y(_04633_)
  );
  XOR2X1 _12550_ (
    .A(_05631_),
    .B(_04632_),
    .Y(_04634_)
  );
  INVX1 _12551_ (
    .A(_04634_),
    .Y(_04635_)
  );
  AOI21X1 _12552_ (
    .A(_05634_),
    .B(_05898_),
    .C(_05633_),
    .Y(_04636_)
  );
  XNOR2X1 _12553_ (
    .A(_04634_),
    .B(_04636_),
    .Y(_04637_)
  );
  NAND2X1 _12554_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05943_),
    .Y(_04638_)
  );
  OAI21X1 _12555_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04637_),
    .C(_04638_),
    .Y(_04639_)
  );
  NOR2X1 _12556_ (
    .A(_05316_),
    .B(_04639_),
    .Y(_04640_)
  );
  NAND2X1 _12557_ (
    .A(_05316_),
    .B(_04639_),
    .Y(_04641_)
  );
  XNOR2X1 _12558_ (
    .A(_05316_),
    .B(_04639_),
    .Y(_04642_)
  );
  XOR2X1 _12559_ (
    .A(_05990_),
    .B(_04642_),
    .Y(_04643_)
  );
  AOI21X1 _12560_ (
    .A(_05361_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04644_)
  );
  OAI21X1 _12561_ (
    .A(_05415_),
    .B(_04643_),
    .C(_04644_),
    .Y(_04645_)
  );
  OAI21X1 _12562_ (
    .A( multiplier_0.reslo_15_ ),
    .B(_05417_),
    .C(_04645_),
    .Y(_04646_)
  );
  INVX1 _12563_ (
    .A(_04646_),
    .Y(_04569_)
  );
  NAND2X1 _12564_ (
    .A(_05904_),
    .B(_05988_),
    .Y(_04647_)
  );
  NAND2X1 _12565_ (
    .A(_05989_),
    .B(_04647_),
    .Y(_04648_)
  );
  AOI21X1 _12566_ (
    .A(_05364_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04649_)
  );
  OAI21X1 _12567_ (
    .A(_05415_),
    .B(_04648_),
    .C(_04649_),
    .Y(_04650_)
  );
  OAI21X1 _12568_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_05417_),
    .C(_04650_),
    .Y(_04651_)
  );
  INVX1 _12569_ (
    .A(_04651_),
    .Y(_04568_)
  );
  XNOR2X1 _12570_ (
    .A(_05910_),
    .B(_05987_),
    .Y(_04652_)
  );
  AOI21X1 _12571_ (
    .A(_05367_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04653_)
  );
  OAI21X1 _12572_ (
    .A(_05415_),
    .B(_04652_),
    .C(_04653_),
    .Y(_04654_)
  );
  OAI21X1 _12573_ (
    .A( multiplier_0.reslo_13_ ),
    .B(_05417_),
    .C(_04654_),
    .Y(_04655_)
  );
  INVX1 _12574_ (
    .A(_04655_),
    .Y(_04567_)
  );
  XNOR2X1 _12575_ (
    .A(_05915_),
    .B(_05986_),
    .Y(_04656_)
  );
  AOI21X1 _12576_ (
    .A(_05370_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04657_)
  );
  OAI21X1 _12577_ (
    .A(_05415_),
    .B(_04656_),
    .C(_04657_),
    .Y(_04658_)
  );
  OAI21X1 _12578_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_05417_),
    .C(_04658_),
    .Y(_04659_)
  );
  INVX1 _12579_ (
    .A(_04659_),
    .Y(_04566_)
  );
  XOR2X1 _12580_ (
    .A(_05923_),
    .B(_05985_),
    .Y(_04660_)
  );
  AOI21X1 _12581_ (
    .A(_05373_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04661_)
  );
  OAI21X1 _12582_ (
    .A(_05415_),
    .B(_04660_),
    .C(_04661_),
    .Y(_04662_)
  );
  OAI21X1 _12583_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_05417_),
    .C(_04662_),
    .Y(_04663_)
  );
  INVX1 _12584_ (
    .A(_04663_),
    .Y(_04565_)
  );
  XNOR2X1 _12585_ (
    .A(_05930_),
    .B(_05984_),
    .Y(_04664_)
  );
  AOI21X1 _12586_ (
    .A(_05376_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04665_)
  );
  OAI21X1 _12587_ (
    .A(_05415_),
    .B(_04664_),
    .C(_04665_),
    .Y(_04666_)
  );
  OAI21X1 _12588_ (
    .A( multiplier_0.reslo_10_ ),
    .B(_05417_),
    .C(_04666_),
    .Y(_04667_)
  );
  INVX1 _12589_ (
    .A(_04667_),
    .Y(_04564_)
  );
  XOR2X1 _12590_ (
    .A(_05938_),
    .B(_05983_),
    .Y(_04668_)
  );
  AOI21X1 _12591_ (
    .A(_05379_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04669_)
  );
  OAI21X1 _12592_ (
    .A(_05415_),
    .B(_04668_),
    .C(_04669_),
    .Y(_04670_)
  );
  OAI21X1 _12593_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_05417_),
    .C(_04670_),
    .Y(_04671_)
  );
  INVX1 _12594_ (
    .A(_04671_),
    .Y(_04563_)
  );
  XNOR2X1 _12595_ (
    .A(_05981_),
    .B(_05982_),
    .Y(_04672_)
  );
  AOI21X1 _12596_ (
    .A(_05382_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04673_)
  );
  OAI21X1 _12597_ (
    .A(_05415_),
    .B(_04672_),
    .C(_04673_),
    .Y(_04674_)
  );
  OAI21X1 _12598_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_05417_),
    .C(_04674_),
    .Y(_04675_)
  );
  INVX1 _12599_ (
    .A(_04675_),
    .Y(_04562_)
  );
  XNOR2X1 _12600_ (
    .A(_05948_),
    .B(_05980_),
    .Y(_04676_)
  );
  INVX1 _12601_ (
    .A(_04676_),
    .Y(_04677_)
  );
  AOI21X1 _12602_ (
    .A(_06288_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04678_)
  );
  OAI21X1 _12603_ (
    .A(_05415_),
    .B(_04677_),
    .C(_04678_),
    .Y(_04679_)
  );
  OAI21X1 _12604_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_05417_),
    .C(_04679_),
    .Y(_04680_)
  );
  INVX1 _12605_ (
    .A(_04680_),
    .Y(_04561_)
  );
  XOR2X1 _12606_ (
    .A(_05952_),
    .B(_05979_),
    .Y(_04681_)
  );
  AOI21X1 _12607_ (
    .A(_06287_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04682_)
  );
  OAI21X1 _12608_ (
    .A(_05415_),
    .B(_04681_),
    .C(_04682_),
    .Y(_04683_)
  );
  OAI21X1 _12609_ (
    .A( multiplier_0.reslo_6_ ),
    .B(_05417_),
    .C(_04683_),
    .Y(_04684_)
  );
  INVX1 _12610_ (
    .A(_04684_),
    .Y(_04560_)
  );
  XNOR2X1 _12611_ (
    .A(_05957_),
    .B(_05978_),
    .Y(_04685_)
  );
  INVX1 _12612_ (
    .A(_04685_),
    .Y(_04686_)
  );
  AOI21X1 _12613_ (
    .A(_06286_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04687_)
  );
  OAI21X1 _12614_ (
    .A(_05415_),
    .B(_04686_),
    .C(_04687_),
    .Y(_04688_)
  );
  OAI21X1 _12615_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_05417_),
    .C(_04688_),
    .Y(_04689_)
  );
  INVX1 _12616_ (
    .A(_04689_),
    .Y(_04559_)
  );
  XOR2X1 _12617_ (
    .A(_05975_),
    .B(_05976_),
    .Y(_04690_)
  );
  INVX1 _12618_ (
    .A(_04690_),
    .Y(_04691_)
  );
  AOI21X1 _12619_ (
    .A(_06285_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04692_)
  );
  OAI21X1 _12620_ (
    .A(_05415_),
    .B(_04691_),
    .C(_04692_),
    .Y(_04693_)
  );
  OAI21X1 _12621_ (
    .A( multiplier_0.reslo_4_ ),
    .B(_05417_),
    .C(_04693_),
    .Y(_04694_)
  );
  INVX1 _12622_ (
    .A(_04694_),
    .Y(_04558_)
  );
  XNOR2X1 _12623_ (
    .A(_05963_),
    .B(_05974_),
    .Y(_04695_)
  );
  INVX1 _12624_ (
    .A(_04695_),
    .Y(_04696_)
  );
  AOI21X1 _12625_ (
    .A(_06284_),
    .B(_05414_),
    .C(_05416_),
    .Y(_04697_)
  );
  OAI21X1 _12626_ (
    .A(_05415_),
    .B(_04696_),
    .C(_04697_),
    .Y(_04698_)
  );
  OAI21X1 _12627_ (
    .A( multiplier_0.reslo_3_ ),
    .B(_05417_),
    .C(_04698_),
    .Y(_04699_)
  );
  INVX1 _12628_ (
    .A(_04699_),
    .Y(_04557_)
  );
  XNOR2X1 _12629_ (
    .A(_05966_),
    .B(_05973_),
    .Y(_04700_)
  );
  NAND2X1 _12630_ (
    .A(_06283_),
    .B(_05414_),
    .Y(_04701_)
  );
  OAI21X1 _12631_ (
    .A(_05415_),
    .B(_04700_),
    .C(_04701_),
    .Y(_04702_)
  );
  OAI21X1 _12632_ (
    .A(_05412_),
    .B(_05415_),
    .C(_04702_),
    .Y(_04703_)
  );
  OAI21X1 _12633_ (
    .A(_05319_),
    .B(_05417_),
    .C(_04703_),
    .Y(_04556_)
  );
  XNOR2X1 _12634_ (
    .A(_05969_),
    .B(_05972_),
    .Y(_04704_)
  );
  NOR2X1 _12635_ (
    .A(_05415_),
    .B(_04704_),
    .Y(_04705_)
  );
  AOI21X1 _12636_ (
    .A(_06282_),
    .B(_05414_),
    .C(_04705_),
    .Y(_04706_)
  );
  NAND2X1 _12637_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_05416_),
    .Y(_04707_)
  );
  OAI21X1 _12638_ (
    .A(_05416_),
    .B(_04706_),
    .C(_04707_),
    .Y(_04555_)
  );
  NAND2X1 _12639_ (
    .A(_05320_),
    .B(_05874_),
    .Y(_04708_)
  );
  NAND2X1 _12640_ (
    .A(_05970_),
    .B(_04708_),
    .Y(_04709_)
  );
  NAND2X1 _12641_ (
    .A(_06275_),
    .B(_05414_),
    .Y(_04710_)
  );
  OAI21X1 _12642_ (
    .A(_05415_),
    .B(_04709_),
    .C(_04710_),
    .Y(_04711_)
  );
  OAI21X1 _12643_ (
    .A(_05412_),
    .B(_05415_),
    .C(_04711_),
    .Y(_04712_)
  );
  OAI21X1 _12644_ (
    .A(_05320_),
    .B(_05417_),
    .C(_04712_),
    .Y(_04554_)
  );
  NAND2X1 _12645_ (
    .A(_06267_),
    .B(_06266_),
    .Y(_04713_)
  );
  OR2X1 _12646_ (
    .A(_06262_),
    .B(_04713_),
    .Y(_04714_)
  );
  NOR2X1 _12647_ (
    .A(_05351_),
    .B(_04714_),
    .Y(_04715_)
  );
  OAI22X1 _12648_ (
    .A( multiplier_0.acc_sel ),
    .B(_05394_),
    .C(_04714_),
    .D(_05358_),
    .Y(_04716_)
  );
  NOR2X1 _12649_ (
    .A(_05412_),
    .B(_04716_),
    .Y(_04717_)
  );
  OR2X1 _12650_ (
    .A(_05412_),
    .B(_04716_),
    .Y(_04718_)
  );
  NOR2X1 _12651_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05485_),
    .Y(_04719_)
  );
  NAND2X1 _12652_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05479_),
    .Y(_04720_)
  );
  NAND2X1 _12653_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05481_),
    .Y(_04721_)
  );
  NAND2X1 _12654_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05481_),
    .Y(_04722_)
  );
  NAND2X1 _12655_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05479_),
    .Y(_04723_)
  );
  OR2X1 _12656_ (
    .A(_04720_),
    .B(_04721_),
    .Y(_04724_)
  );
  NAND2X1 _12657_ (
    .A(_04720_),
    .B(_04721_),
    .Y(_04725_)
  );
  OAI21X1 _12658_ (
    .A(_04722_),
    .B(_04723_),
    .C(_04725_),
    .Y(_04726_)
  );
  NAND3X1 _12659_ (
    .A(_04719_),
    .B(_04724_),
    .C(_04725_),
    .Y(_04727_)
  );
  OAI21X1 _12660_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05485_),
    .C(_04726_),
    .Y(_04728_)
  );
  NAND2X1 _12661_ (
    .A(_04727_),
    .B(_04728_),
    .Y(_04729_)
  );
  NOR2X1 _12662_ (
    .A(_05298_),
    .B(_05332_),
    .Y(_04730_)
  );
  NAND2X1 _12663_ (
    .A( multiplier_0.op1_15_ ),
    .B( multiplier_0.sign_sel ),
    .Y(_04731_)
  );
  AND2X1 _12664_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05450_),
    .Y(_04732_)
  );
  NAND3X1 _12665_ (
    .A(_05447_),
    .B(_05450_),
    .C(_04730_),
    .Y(_04733_)
  );
  INVX1 _12666_ (
    .A(_04733_),
    .Y(_04734_)
  );
  NAND2X1 _12667_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05444_),
    .Y(_04735_)
  );
  AOI22X1 _12668_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05447_),
    .C(_05450_),
    .D(_04730_),
    .Y(_04736_)
  );
  OR2X1 _12669_ (
    .A(_04734_),
    .B(_04736_),
    .Y(_04737_)
  );
  NOR2X1 _12670_ (
    .A(_04735_),
    .B(_04737_),
    .Y(_04738_)
  );
  NOR2X1 _12671_ (
    .A(_04734_),
    .B(_04738_),
    .Y(_04739_)
  );
  NOR2X1 _12672_ (
    .A(_04729_),
    .B(_04739_),
    .Y(_04740_)
  );
  NAND2X1 _12673_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05479_),
    .Y(_04741_)
  );
  OR2X1 _12674_ (
    .A(_04722_),
    .B(_04741_),
    .Y(_04742_)
  );
  NOR2X1 _12675_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05485_),
    .Y(_04743_)
  );
  NAND2X1 _12676_ (
    .A(_04722_),
    .B(_04741_),
    .Y(_04744_)
  );
  NAND2X1 _12677_ (
    .A(_04742_),
    .B(_04744_),
    .Y(_04745_)
  );
  NAND3X1 _12678_ (
    .A(_04742_),
    .B(_04743_),
    .C(_04744_),
    .Y(_04746_)
  );
  OAI21X1 _12679_ (
    .A(_04722_),
    .B(_04741_),
    .C(_04746_),
    .Y(_04747_)
  );
  NAND2X1 _12680_ (
    .A(_04729_),
    .B(_04739_),
    .Y(_04748_)
  );
  XNOR2X1 _12681_ (
    .A(_04729_),
    .B(_04739_),
    .Y(_04749_)
  );
  AOI21X1 _12682_ (
    .A(_04747_),
    .B(_04748_),
    .C(_04740_),
    .Y(_04750_)
  );
  NAND2X1 _12683_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05429_),
    .Y(_04751_)
  );
  NAND2X1 _12684_ (
    .A(_05429_),
    .B(_04730_),
    .Y(_04752_)
  );
  INVX1 _12685_ (
    .A(_04752_),
    .Y(_04753_)
  );
  NOR2X1 _12686_ (
    .A(_05422_),
    .B(_04731_),
    .Y(_04754_)
  );
  NAND2X1 _12687_ (
    .A(_05420_),
    .B(_04754_),
    .Y(_04755_)
  );
  OR2X1 _12688_ (
    .A(_04752_),
    .B(_04755_),
    .Y(_04756_)
  );
  XNOR2X1 _12689_ (
    .A(_04735_),
    .B(_04737_),
    .Y(_04757_)
  );
  AOI21X1 _12690_ (
    .A(_05419_),
    .B(_05422_),
    .C(_04731_),
    .Y(_04758_)
  );
  OAI21X1 _12691_ (
    .A(_04753_),
    .B(_04758_),
    .C(_04756_),
    .Y(_04759_)
  );
  OR2X1 _12692_ (
    .A(_04757_),
    .B(_04759_),
    .Y(_04760_)
  );
  NAND2X1 _12693_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05444_),
    .Y(_04761_)
  );
  OAI21X1 _12694_ (
    .A(_05447_),
    .B(_05450_),
    .C(_04730_),
    .Y(_04762_)
  );
  NOR2X1 _12695_ (
    .A(_04734_),
    .B(_04762_),
    .Y(_04763_)
  );
  NAND3X1 _12696_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05444_),
    .C(_04763_),
    .Y(_04764_)
  );
  INVX1 _12697_ (
    .A(_04764_),
    .Y(_04765_)
  );
  OAI21X1 _12698_ (
    .A(_04734_),
    .B(_04762_),
    .C(_04761_),
    .Y(_04766_)
  );
  NAND2X1 _12699_ (
    .A(_04764_),
    .B(_04766_),
    .Y(_04767_)
  );
  XNOR2X1 _12700_ (
    .A(_04759_),
    .B(_04767_),
    .Y(_04768_)
  );
  AOI21X1 _12701_ (
    .A(_04756_),
    .B(_04760_),
    .C(_04768_),
    .Y(_04769_)
  );
  INVX1 _12702_ (
    .A(_04769_),
    .Y(_04770_)
  );
  XOR2X1 _12703_ (
    .A(_04747_),
    .B(_04749_),
    .Y(_04771_)
  );
  NAND3X1 _12704_ (
    .A(_04756_),
    .B(_04760_),
    .C(_04768_),
    .Y(_04772_)
  );
  NAND2X1 _12705_ (
    .A(_04770_),
    .B(_04772_),
    .Y(_04773_)
  );
  OAI21X1 _12706_ (
    .A(_04771_),
    .B(_04773_),
    .C(_04770_),
    .Y(_04774_)
  );
  OAI21X1 _12707_ (
    .A(_04722_),
    .B(_04723_),
    .C(_04727_),
    .Y(_04775_)
  );
  NOR2X1 _12708_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05485_),
    .Y(_04776_)
  );
  NAND2X1 _12709_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05481_),
    .Y(_04777_)
  );
  NAND2X1 _12710_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05479_),
    .Y(_04778_)
  );
  XOR2X1 _12711_ (
    .A(_04723_),
    .B(_04777_),
    .Y(_04779_)
  );
  NAND2X1 _12712_ (
    .A(_04776_),
    .B(_04779_),
    .Y(_04780_)
  );
  XNOR2X1 _12713_ (
    .A(_04776_),
    .B(_04779_),
    .Y(_04781_)
  );
  NOR2X1 _12714_ (
    .A(_04734_),
    .B(_04765_),
    .Y(_04782_)
  );
  OAI21X1 _12715_ (
    .A(_04761_),
    .B(_04762_),
    .C(_04733_),
    .Y(_04783_)
  );
  NOR2X1 _12716_ (
    .A(_04781_),
    .B(_04782_),
    .Y(_04784_)
  );
  XOR2X1 _12717_ (
    .A(_04781_),
    .B(_04783_),
    .Y(_04785_)
  );
  AOI21X1 _12718_ (
    .A(_04724_),
    .B(_04727_),
    .C(_04785_),
    .Y(_04786_)
  );
  XOR2X1 _12719_ (
    .A(_04775_),
    .B(_04785_),
    .Y(_04787_)
  );
  AOI21X1 _12720_ (
    .A(_05444_),
    .B(_04730_),
    .C(_04763_),
    .Y(_04788_)
  );
  OAI21X1 _12721_ (
    .A(_04765_),
    .B(_04788_),
    .C(_04759_),
    .Y(_04789_)
  );
  INVX1 _12722_ (
    .A(_04789_),
    .Y(_04790_)
  );
  NOR2X1 _12723_ (
    .A(_04756_),
    .B(_04790_),
    .Y(_04791_)
  );
  INVX1 _12724_ (
    .A(_04791_),
    .Y(_04792_)
  );
  XNOR2X1 _12725_ (
    .A(_04756_),
    .B(_04789_),
    .Y(_04793_)
  );
  INVX1 _12726_ (
    .A(_04793_),
    .Y(_04794_)
  );
  XNOR2X1 _12727_ (
    .A(_04787_),
    .B(_04793_),
    .Y(_04795_)
  );
  NAND2X1 _12728_ (
    .A(_04774_),
    .B(_04795_),
    .Y(_04796_)
  );
  XNOR2X1 _12729_ (
    .A(_04774_),
    .B(_04795_),
    .Y(_04797_)
  );
  XOR2X1 _12730_ (
    .A(_04750_),
    .B(_04797_),
    .Y(_04798_)
  );
  NAND2X1 _12731_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05444_),
    .Y(_04799_)
  );
  NAND2X1 _12732_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05447_),
    .Y(_04800_)
  );
  NAND2X1 _12733_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05450_),
    .Y(_04801_)
  );
  NAND3X1 _12734_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05447_),
    .C(_04732_),
    .Y(_04802_)
  );
  XOR2X1 _12735_ (
    .A(_04732_),
    .B(_04800_),
    .Y(_04803_)
  );
  XNOR2X1 _12736_ (
    .A(_04799_),
    .B(_04803_),
    .Y(_04804_)
  );
  OAI21X1 _12737_ (
    .A(_04759_),
    .B(_04804_),
    .C(_04756_),
    .Y(_04805_)
  );
  XOR2X1 _12738_ (
    .A(_04757_),
    .B(_04759_),
    .Y(_04806_)
  );
  NAND2X1 _12739_ (
    .A(_04805_),
    .B(_04806_),
    .Y(_04807_)
  );
  NAND2X1 _12740_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05479_),
    .Y(_04808_)
  );
  NAND2X1 _12741_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05481_),
    .Y(_04809_)
  );
  NOR2X1 _12742_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05485_),
    .Y(_04810_)
  );
  INVX1 _12743_ (
    .A(_04810_),
    .Y(_04811_)
  );
  OAI21X1 _12744_ (
    .A(_05299_),
    .B(_05482_),
    .C(_04808_),
    .Y(_04812_)
  );
  OAI21X1 _12745_ (
    .A(_04741_),
    .B(_04809_),
    .C(_04812_),
    .Y(_04813_)
  );
  OAI22X1 _12746_ (
    .A(_04741_),
    .B(_04809_),
    .C(_04811_),
    .D(_04813_),
    .Y(_04814_)
  );
  OAI21X1 _12747_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05485_),
    .C(_04745_),
    .Y(_04815_)
  );
  NAND2X1 _12748_ (
    .A(_04746_),
    .B(_04815_),
    .Y(_04816_)
  );
  OAI21X1 _12749_ (
    .A(_04799_),
    .B(_04803_),
    .C(_04802_),
    .Y(_04817_)
  );
  INVX1 _12750_ (
    .A(_04817_),
    .Y(_04818_)
  );
  XNOR2X1 _12751_ (
    .A(_04816_),
    .B(_04818_),
    .Y(_04819_)
  );
  INVX1 _12752_ (
    .A(_04819_),
    .Y(_04820_)
  );
  NAND2X1 _12753_ (
    .A(_04814_),
    .B(_04820_),
    .Y(_04821_)
  );
  XOR2X1 _12754_ (
    .A(_04814_),
    .B(_04819_),
    .Y(_04822_)
  );
  XNOR2X1 _12755_ (
    .A(_04805_),
    .B(_04806_),
    .Y(_04823_)
  );
  OAI21X1 _12756_ (
    .A(_04822_),
    .B(_04823_),
    .C(_04807_),
    .Y(_04824_)
  );
  XOR2X1 _12757_ (
    .A(_04771_),
    .B(_04773_),
    .Y(_04825_)
  );
  NAND2X1 _12758_ (
    .A(_04824_),
    .B(_04825_),
    .Y(_04826_)
  );
  OAI21X1 _12759_ (
    .A(_04816_),
    .B(_04818_),
    .C(_04821_),
    .Y(_04827_)
  );
  INVX1 _12760_ (
    .A(_04827_),
    .Y(_04828_)
  );
  XNOR2X1 _12761_ (
    .A(_04824_),
    .B(_04825_),
    .Y(_04829_)
  );
  OAI21X1 _12762_ (
    .A(_04828_),
    .B(_04829_),
    .C(_04826_),
    .Y(_04830_)
  );
  NAND2X1 _12763_ (
    .A(_04798_),
    .B(_04830_),
    .Y(_04831_)
  );
  XOR2X1 _12764_ (
    .A(_04798_),
    .B(_04830_),
    .Y(_04832_)
  );
  XNOR2X1 _12765_ (
    .A(_04827_),
    .B(_04829_),
    .Y(_04833_)
  );
  NAND2X1 _12766_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05429_),
    .Y(_04834_)
  );
  OAI21X1 _12767_ (
    .A(_04617_),
    .B(_04754_),
    .C(_04755_),
    .Y(_04835_)
  );
  OAI21X1 _12768_ (
    .A(_04834_),
    .B(_04835_),
    .C(_04755_),
    .Y(_04836_)
  );
  NAND2X1 _12769_ (
    .A(_04755_),
    .B(_04758_),
    .Y(_04837_)
  );
  NAND2X1 _12770_ (
    .A(_04751_),
    .B(_04837_),
    .Y(_04838_)
  );
  OAI21X1 _12771_ (
    .A(_04752_),
    .B(_04837_),
    .C(_04838_),
    .Y(_04839_)
  );
  INVX1 _12772_ (
    .A(_04839_),
    .Y(_04840_)
  );
  NAND2X1 _12773_ (
    .A(_04836_),
    .B(_04840_),
    .Y(_04841_)
  );
  NAND2X1 _12774_ (
    .A( multiplier_0.op1_12_ ),
    .B(_05444_),
    .Y(_04842_)
  );
  NAND2X1 _12775_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05447_),
    .Y(_04843_)
  );
  NAND2X1 _12776_ (
    .A( multiplier_0.op1_13_ ),
    .B(_05450_),
    .Y(_04844_)
  );
  XNOR2X1 _12777_ (
    .A(_04801_),
    .B(_04843_),
    .Y(_04845_)
  );
  XOR2X1 _12778_ (
    .A(_04842_),
    .B(_04845_),
    .Y(_04846_)
  );
  XNOR2X1 _12779_ (
    .A(_04836_),
    .B(_04839_),
    .Y(_04847_)
  );
  NAND2X1 _12780_ (
    .A(_04846_),
    .B(_04847_),
    .Y(_04848_)
  );
  XNOR2X1 _12781_ (
    .A(_04759_),
    .B(_04804_),
    .Y(_04849_)
  );
  AOI21X1 _12782_ (
    .A(_04841_),
    .B(_04848_),
    .C(_04849_),
    .Y(_04850_)
  );
  INVX1 _12783_ (
    .A(_04850_),
    .Y(_04851_)
  );
  NAND2X1 _12784_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05479_),
    .Y(_04852_)
  );
  NAND2X1 _12785_ (
    .A( multiplier_0.op1_10_ ),
    .B(_05481_),
    .Y(_04853_)
  );
  NOR2X1 _12786_ (
    .A( multiplier_0.op1_9_ ),
    .B(_05485_),
    .Y(_04854_)
  );
  INVX1 _12787_ (
    .A(_04854_),
    .Y(_04855_)
  );
  NAND2X1 _12788_ (
    .A(_04809_),
    .B(_04852_),
    .Y(_04856_)
  );
  OAI21X1 _12789_ (
    .A(_04808_),
    .B(_04853_),
    .C(_04856_),
    .Y(_04857_)
  );
  OAI22X1 _12790_ (
    .A(_04808_),
    .B(_04853_),
    .C(_04855_),
    .D(_04857_),
    .Y(_04858_)
  );
  XNOR2X1 _12791_ (
    .A(_04811_),
    .B(_04813_),
    .Y(_04859_)
  );
  OAI22X1 _12792_ (
    .A(_04800_),
    .B(_04844_),
    .C(_04845_),
    .D(_04842_),
    .Y(_04860_)
  );
  INVX1 _12793_ (
    .A(_04860_),
    .Y(_04861_)
  );
  XOR2X1 _12794_ (
    .A(_04859_),
    .B(_04860_),
    .Y(_04862_)
  );
  INVX1 _12795_ (
    .A(_04862_),
    .Y(_04863_)
  );
  NAND2X1 _12796_ (
    .A(_04858_),
    .B(_04863_),
    .Y(_04864_)
  );
  XOR2X1 _12797_ (
    .A(_04858_),
    .B(_04862_),
    .Y(_04865_)
  );
  NAND3X1 _12798_ (
    .A(_04841_),
    .B(_04848_),
    .C(_04849_),
    .Y(_04866_)
  );
  NAND2X1 _12799_ (
    .A(_04851_),
    .B(_04866_),
    .Y(_04867_)
  );
  OAI21X1 _12800_ (
    .A(_04865_),
    .B(_04867_),
    .C(_04851_),
    .Y(_04868_)
  );
  XOR2X1 _12801_ (
    .A(_04822_),
    .B(_04823_),
    .Y(_04869_)
  );
  NAND2X1 _12802_ (
    .A(_04868_),
    .B(_04869_),
    .Y(_04870_)
  );
  OAI21X1 _12803_ (
    .A(_04859_),
    .B(_04861_),
    .C(_04864_),
    .Y(_04871_)
  );
  INVX1 _12804_ (
    .A(_04871_),
    .Y(_04872_)
  );
  XNOR2X1 _12805_ (
    .A(_04868_),
    .B(_04869_),
    .Y(_04873_)
  );
  OAI21X1 _12806_ (
    .A(_04872_),
    .B(_04873_),
    .C(_04870_),
    .Y(_04874_)
  );
  NAND2X1 _12807_ (
    .A(_04833_),
    .B(_04874_),
    .Y(_04875_)
  );
  NAND3X1 _12808_ (
    .A(_04832_),
    .B(_04833_),
    .C(_04874_),
    .Y(_04876_)
  );
  XNOR2X1 _12809_ (
    .A(_04832_),
    .B(_04875_),
    .Y(_04877_)
  );
  INVX1 _12810_ (
    .A(_04877_),
    .Y(_04878_)
  );
  XNOR2X1 _12811_ (
    .A(_04833_),
    .B(_04874_),
    .Y(_04879_)
  );
  XNOR2X1 _12812_ (
    .A(_04871_),
    .B(_04873_),
    .Y(_04880_)
  );
  OAI22X1 _12813_ (
    .A(_05616_),
    .B(_04616_),
    .C(_04619_),
    .D(_04615_),
    .Y(_04881_)
  );
  XNOR2X1 _12814_ (
    .A(_04834_),
    .B(_04835_),
    .Y(_04882_)
  );
  INVX1 _12815_ (
    .A(_04882_),
    .Y(_04883_)
  );
  NAND2X1 _12816_ (
    .A(_04881_),
    .B(_04883_),
    .Y(_04884_)
  );
  NAND2X1 _12817_ (
    .A( multiplier_0.op1_11_ ),
    .B(_05444_),
    .Y(_04885_)
  );
  XNOR2X1 _12818_ (
    .A(_04610_),
    .B(_04844_),
    .Y(_04886_)
  );
  XNOR2X1 _12819_ (
    .A(_04885_),
    .B(_04886_),
    .Y(_04887_)
  );
  XOR2X1 _12820_ (
    .A(_04881_),
    .B(_04882_),
    .Y(_04888_)
  );
  OAI21X1 _12821_ (
    .A(_04887_),
    .B(_04888_),
    .C(_04884_),
    .Y(_04889_)
  );
  XOR2X1 _12822_ (
    .A(_04846_),
    .B(_04847_),
    .Y(_04890_)
  );
  NAND2X1 _12823_ (
    .A(_04889_),
    .B(_04890_),
    .Y(_04891_)
  );
  NOR2X1 _12824_ (
    .A( multiplier_0.op1_8_ ),
    .B(_05485_),
    .Y(_04892_)
  );
  INVX1 _12825_ (
    .A(_04892_),
    .Y(_04893_)
  );
  NAND2X1 _12826_ (
    .A(_05999_),
    .B(_04853_),
    .Y(_04894_)
  );
  OAI21X1 _12827_ (
    .A(_05998_),
    .B(_04852_),
    .C(_04894_),
    .Y(_04895_)
  );
  OAI22X1 _12828_ (
    .A(_05998_),
    .B(_04852_),
    .C(_04893_),
    .D(_04895_),
    .Y(_04896_)
  );
  XNOR2X1 _12829_ (
    .A(_04855_),
    .B(_04857_),
    .Y(_04897_)
  );
  OAI22X1 _12830_ (
    .A(_04609_),
    .B(_04843_),
    .C(_04885_),
    .D(_04886_),
    .Y(_04898_)
  );
  INVX1 _12831_ (
    .A(_04898_),
    .Y(_04899_)
  );
  XNOR2X1 _12832_ (
    .A(_04897_),
    .B(_04899_),
    .Y(_04900_)
  );
  INVX1 _12833_ (
    .A(_04900_),
    .Y(_04901_)
  );
  NAND2X1 _12834_ (
    .A(_04896_),
    .B(_04901_),
    .Y(_04902_)
  );
  XOR2X1 _12835_ (
    .A(_04896_),
    .B(_04900_),
    .Y(_04903_)
  );
  XNOR2X1 _12836_ (
    .A(_04889_),
    .B(_04890_),
    .Y(_04904_)
  );
  OAI21X1 _12837_ (
    .A(_04903_),
    .B(_04904_),
    .C(_04891_),
    .Y(_04905_)
  );
  XOR2X1 _12838_ (
    .A(_04865_),
    .B(_04867_),
    .Y(_04906_)
  );
  NAND2X1 _12839_ (
    .A(_04905_),
    .B(_04906_),
    .Y(_04907_)
  );
  OAI21X1 _12840_ (
    .A(_04897_),
    .B(_04899_),
    .C(_04902_),
    .Y(_04908_)
  );
  INVX1 _12841_ (
    .A(_04908_),
    .Y(_04909_)
  );
  XNOR2X1 _12842_ (
    .A(_04905_),
    .B(_04906_),
    .Y(_04910_)
  );
  OAI21X1 _12843_ (
    .A(_04909_),
    .B(_04910_),
    .C(_04907_),
    .Y(_04911_)
  );
  NAND2X1 _12844_ (
    .A(_04880_),
    .B(_04911_),
    .Y(_04912_)
  );
  NOR2X1 _12845_ (
    .A(_04879_),
    .B(_04912_),
    .Y(_04913_)
  );
  XOR2X1 _12846_ (
    .A(_04879_),
    .B(_04912_),
    .Y(_04914_)
  );
  XNOR2X1 _12847_ (
    .A(_04880_),
    .B(_04911_),
    .Y(_04915_)
  );
  XNOR2X1 _12848_ (
    .A(_04908_),
    .B(_04910_),
    .Y(_04916_)
  );
  OAI21X1 _12849_ (
    .A(_04613_),
    .B(_04623_),
    .C(_04622_),
    .Y(_04917_)
  );
  XOR2X1 _12850_ (
    .A(_04887_),
    .B(_04888_),
    .Y(_04918_)
  );
  NAND2X1 _12851_ (
    .A(_04917_),
    .B(_04918_),
    .Y(_04919_)
  );
  OAI22X1 _12852_ (
    .A(_05596_),
    .B(_05999_),
    .C(_06001_),
    .D(_05997_),
    .Y(_04920_)
  );
  XNOR2X1 _12853_ (
    .A(_04893_),
    .B(_04895_),
    .Y(_04921_)
  );
  OAI21X1 _12854_ (
    .A(_04608_),
    .B(_04612_),
    .C(_04611_),
    .Y(_04922_)
  );
  INVX1 _12855_ (
    .A(_04922_),
    .Y(_04923_)
  );
  XNOR2X1 _12856_ (
    .A(_04921_),
    .B(_04923_),
    .Y(_04924_)
  );
  INVX1 _12857_ (
    .A(_04924_),
    .Y(_04925_)
  );
  NAND2X1 _12858_ (
    .A(_04920_),
    .B(_04925_),
    .Y(_04926_)
  );
  XOR2X1 _12859_ (
    .A(_04920_),
    .B(_04924_),
    .Y(_04927_)
  );
  XNOR2X1 _12860_ (
    .A(_04917_),
    .B(_04918_),
    .Y(_04928_)
  );
  OAI21X1 _12861_ (
    .A(_04927_),
    .B(_04928_),
    .C(_04919_),
    .Y(_04929_)
  );
  XOR2X1 _12862_ (
    .A(_04903_),
    .B(_04904_),
    .Y(_04930_)
  );
  NAND2X1 _12863_ (
    .A(_04929_),
    .B(_04930_),
    .Y(_04931_)
  );
  OAI21X1 _12864_ (
    .A(_04921_),
    .B(_04923_),
    .C(_04926_),
    .Y(_04932_)
  );
  INVX1 _12865_ (
    .A(_04932_),
    .Y(_04933_)
  );
  XNOR2X1 _12866_ (
    .A(_04929_),
    .B(_04930_),
    .Y(_04934_)
  );
  OAI21X1 _12867_ (
    .A(_04933_),
    .B(_04934_),
    .C(_04931_),
    .Y(_04935_)
  );
  NAND2X1 _12868_ (
    .A(_04916_),
    .B(_04935_),
    .Y(_04936_)
  );
  OR2X1 _12869_ (
    .A(_04915_),
    .B(_04936_),
    .Y(_04937_)
  );
  XOR2X1 _12870_ (
    .A(_04915_),
    .B(_04936_),
    .Y(_04938_)
  );
  INVX1 _12871_ (
    .A(_04938_),
    .Y(_04939_)
  );
  XNOR2X1 _12872_ (
    .A(_04916_),
    .B(_04935_),
    .Y(_04940_)
  );
  XNOR2X1 _12873_ (
    .A(_04932_),
    .B(_04934_),
    .Y(_04941_)
  );
  OAI21X1 _12874_ (
    .A(_04606_),
    .B(_04626_),
    .C(_04625_),
    .Y(_04942_)
  );
  XOR2X1 _12875_ (
    .A(_04927_),
    .B(_04928_),
    .Y(_04943_)
  );
  NAND2X1 _12876_ (
    .A(_04942_),
    .B(_04943_),
    .Y(_04944_)
  );
  OAI21X1 _12877_ (
    .A(_06002_),
    .B(_04602_),
    .C(_04605_),
    .Y(_04945_)
  );
  INVX1 _12878_ (
    .A(_04945_),
    .Y(_04946_)
  );
  XNOR2X1 _12879_ (
    .A(_04942_),
    .B(_04943_),
    .Y(_04947_)
  );
  OAI21X1 _12880_ (
    .A(_04946_),
    .B(_04947_),
    .C(_04944_),
    .Y(_04948_)
  );
  NAND2X1 _12881_ (
    .A(_04941_),
    .B(_04948_),
    .Y(_04949_)
  );
  NOR2X1 _12882_ (
    .A(_04940_),
    .B(_04949_),
    .Y(_04950_)
  );
  XOR2X1 _12883_ (
    .A(_04940_),
    .B(_04949_),
    .Y(_04951_)
  );
  OAI21X1 _12884_ (
    .A(_05993_),
    .B(_04629_),
    .C(_04628_),
    .Y(_04952_)
  );
  XNOR2X1 _12885_ (
    .A(_04945_),
    .B(_04947_),
    .Y(_04953_)
  );
  NAND2X1 _12886_ (
    .A(_04952_),
    .B(_04953_),
    .Y(_04954_)
  );
  XNOR2X1 _12887_ (
    .A(_04941_),
    .B(_04948_),
    .Y(_04955_)
  );
  OR2X1 _12888_ (
    .A(_04954_),
    .B(_04955_),
    .Y(_04956_)
  );
  XOR2X1 _12889_ (
    .A(_04954_),
    .B(_04955_),
    .Y(_04957_)
  );
  INVX1 _12890_ (
    .A(_04957_),
    .Y(_04958_)
  );
  XNOR2X1 _12891_ (
    .A(_04952_),
    .B(_04953_),
    .Y(_04959_)
  );
  NOR2X1 _12892_ (
    .A(_04631_),
    .B(_04959_),
    .Y(_04960_)
  );
  OAI21X1 _12893_ (
    .A(_04635_),
    .B(_04636_),
    .C(_04633_),
    .Y(_04961_)
  );
  XOR2X1 _12894_ (
    .A(_04631_),
    .B(_04959_),
    .Y(_04962_)
  );
  AOI21X1 _12895_ (
    .A(_04961_),
    .B(_04962_),
    .C(_04960_),
    .Y(_04963_)
  );
  OAI21X1 _12896_ (
    .A(_04958_),
    .B(_04963_),
    .C(_04956_),
    .Y(_04964_)
  );
  AOI21X1 _12897_ (
    .A(_04951_),
    .B(_04964_),
    .C(_04950_),
    .Y(_04965_)
  );
  OAI21X1 _12898_ (
    .A(_04939_),
    .B(_04965_),
    .C(_04937_),
    .Y(_04966_)
  );
  AOI21X1 _12899_ (
    .A(_04914_),
    .B(_04966_),
    .C(_04913_),
    .Y(_04967_)
  );
  OAI21X1 _12900_ (
    .A(_04878_),
    .B(_04967_),
    .C(_04876_),
    .Y(_04968_)
  );
  OAI21X1 _12901_ (
    .A(_04750_),
    .B(_04797_),
    .C(_04796_),
    .Y(_04969_)
  );
  NOR2X1 _12902_ (
    .A(_04784_),
    .B(_04786_),
    .Y(_04970_)
  );
  OAI21X1 _12903_ (
    .A(_04787_),
    .B(_04794_),
    .C(_04792_),
    .Y(_04971_)
  );
  INVX1 _12904_ (
    .A(_04971_),
    .Y(_04972_)
  );
  OAI21X1 _12905_ (
    .A(_04721_),
    .B(_04778_),
    .C(_04780_),
    .Y(_04973_)
  );
  NOR2X1 _12906_ (
    .A( multiplier_0.op1_14_ ),
    .B(_05485_),
    .Y(_04974_)
  );
  NAND3X1 _12907_ (
    .A(_05479_),
    .B(_05481_),
    .C(_04730_),
    .Y(_04975_)
  );
  INVX1 _12908_ (
    .A(_04975_),
    .Y(_04976_)
  );
  OAI21X1 _12909_ (
    .A(_05482_),
    .B(_04731_),
    .C(_04778_),
    .Y(_04977_)
  );
  NAND2X1 _12910_ (
    .A(_04975_),
    .B(_04977_),
    .Y(_04978_)
  );
  XOR2X1 _12911_ (
    .A(_04974_),
    .B(_04978_),
    .Y(_04979_)
  );
  NOR2X1 _12912_ (
    .A(_04782_),
    .B(_04979_),
    .Y(_04980_)
  );
  NAND2X1 _12913_ (
    .A(_04782_),
    .B(_04979_),
    .Y(_04981_)
  );
  XOR2X1 _12914_ (
    .A(_04783_),
    .B(_04979_),
    .Y(_04982_)
  );
  XOR2X1 _12915_ (
    .A(_04973_),
    .B(_04982_),
    .Y(_04983_)
  );
  XOR2X1 _12916_ (
    .A(_04793_),
    .B(_04983_),
    .Y(_04984_)
  );
  XNOR2X1 _12917_ (
    .A(_04971_),
    .B(_04984_),
    .Y(_04985_)
  );
  OAI21X1 _12918_ (
    .A(_04784_),
    .B(_04786_),
    .C(_04985_),
    .Y(_04986_)
  );
  XNOR2X1 _12919_ (
    .A(_04970_),
    .B(_04985_),
    .Y(_04987_)
  );
  NAND2X1 _12920_ (
    .A(_04969_),
    .B(_04987_),
    .Y(_04988_)
  );
  XNOR2X1 _12921_ (
    .A(_04969_),
    .B(_04987_),
    .Y(_04989_)
  );
  NOR2X1 _12922_ (
    .A(_04831_),
    .B(_04989_),
    .Y(_04990_)
  );
  XOR2X1 _12923_ (
    .A(_04831_),
    .B(_04989_),
    .Y(_04991_)
  );
  XNOR2X1 _12924_ (
    .A(_04968_),
    .B(_04991_),
    .Y(_04992_)
  );
  NAND2X1 _12925_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04992_),
    .Y(_04993_)
  );
  AOI21X1 _12926_ (
    .A(_04968_),
    .B(_04991_),
    .C(_04990_),
    .Y(_04994_)
  );
  OAI21X1 _12927_ (
    .A(_04972_),
    .B(_04984_),
    .C(_04986_),
    .Y(_04995_)
  );
  OAI21X1 _12928_ (
    .A(_04794_),
    .B(_04983_),
    .C(_04792_),
    .Y(_04996_)
  );
  AOI21X1 _12929_ (
    .A(_04973_),
    .B(_04981_),
    .C(_04980_),
    .Y(_04997_)
  );
  AOI21X1 _12930_ (
    .A(_04974_),
    .B(_04977_),
    .C(_04976_),
    .Y(_04998_)
  );
  OAI21X1 _12931_ (
    .A(_05479_),
    .B(_05481_),
    .C(_04730_),
    .Y(_04999_)
  );
  OAI22X1 _12932_ (
    .A( multiplier_0.op1_15_ ),
    .B(_05485_),
    .C(_04976_),
    .D(_04999_),
    .Y(_05000_)
  );
  AOI21X1 _12933_ (
    .A(_04998_),
    .B(_05000_),
    .C(_04976_),
    .Y(_05001_)
  );
  XNOR2X1 _12934_ (
    .A(_04783_),
    .B(_05001_),
    .Y(_05002_)
  );
  XNOR2X1 _12935_ (
    .A(_04793_),
    .B(_05002_),
    .Y(_05003_)
  );
  XNOR2X1 _12936_ (
    .A(_04997_),
    .B(_05003_),
    .Y(_05004_)
  );
  XNOR2X1 _12937_ (
    .A(_04996_),
    .B(_05004_),
    .Y(_05005_)
  );
  XNOR2X1 _12938_ (
    .A(_04995_),
    .B(_05005_),
    .Y(_05006_)
  );
  XNOR2X1 _12939_ (
    .A(_04988_),
    .B(_05006_),
    .Y(_05007_)
  );
  XNOR2X1 _12940_ (
    .A(_04994_),
    .B(_05007_),
    .Y(_05008_)
  );
  OAI21X1 _12941_ (
    .A(_05332_),
    .B(_05008_),
    .C(_05334_),
    .Y(_05009_)
  );
  NAND2X1 _12942_ (
    .A(_04993_),
    .B(_05009_),
    .Y(_05010_)
  );
  NAND3X1 _12943_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_04993_),
    .C(_05009_),
    .Y(_05011_)
  );
  XOR2X1 _12944_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_05010_),
    .Y(_05012_)
  );
  XNOR2X1 _12945_ (
    .A(_04877_),
    .B(_04967_),
    .Y(_05013_)
  );
  OAI21X1 _12946_ (
    .A(_05334_),
    .B(_05013_),
    .C(_05009_),
    .Y(_05014_)
  );
  NAND2X1 _12947_ (
    .A(_05321_),
    .B(_05014_),
    .Y(_05015_)
  );
  OR2X1 _12948_ (
    .A(_05321_),
    .B(_05014_),
    .Y(_05016_)
  );
  INVX1 _12949_ (
    .A(_05016_),
    .Y(_05017_)
  );
  XOR2X1 _12950_ (
    .A(_04914_),
    .B(_04966_),
    .Y(_05018_)
  );
  OAI21X1 _12951_ (
    .A(_05334_),
    .B(_05018_),
    .C(_05009_),
    .Y(_05019_)
  );
  OR2X1 _12952_ (
    .A(_05322_),
    .B(_05019_),
    .Y(_05020_)
  );
  XOR2X1 _12953_ (
    .A( multiplier_0.reshi_12_ ),
    .B(_05019_),
    .Y(_05021_)
  );
  XNOR2X1 _12954_ (
    .A(_04938_),
    .B(_04965_),
    .Y(_05022_)
  );
  OAI21X1 _12955_ (
    .A(_05334_),
    .B(_05022_),
    .C(_05009_),
    .Y(_05023_)
  );
  NAND2X1 _12956_ (
    .A(_05323_),
    .B(_05023_),
    .Y(_05024_)
  );
  OR2X1 _12957_ (
    .A(_05323_),
    .B(_05023_),
    .Y(_05025_)
  );
  INVX1 _12958_ (
    .A(_05025_),
    .Y(_05026_)
  );
  XOR2X1 _12959_ (
    .A(_04951_),
    .B(_04964_),
    .Y(_05027_)
  );
  OR2X1 _12960_ (
    .A(_05334_),
    .B(_05027_),
    .Y(_05028_)
  );
  AND2X1 _12961_ (
    .A(_05009_),
    .B(_05028_),
    .Y(_05029_)
  );
  NAND2X1 _12962_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_05029_),
    .Y(_05030_)
  );
  XNOR2X1 _12963_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_05029_),
    .Y(_05031_)
  );
  XNOR2X1 _12964_ (
    .A(_04958_),
    .B(_04963_),
    .Y(_05032_)
  );
  NAND2X1 _12965_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05032_),
    .Y(_05033_)
  );
  NAND2X1 _12966_ (
    .A(_05009_),
    .B(_05033_),
    .Y(_05034_)
  );
  OR2X1 _12967_ (
    .A(_05324_),
    .B(_05034_),
    .Y(_05035_)
  );
  INVX1 _12968_ (
    .A(_05035_),
    .Y(_05036_)
  );
  NAND2X1 _12969_ (
    .A(_05324_),
    .B(_05034_),
    .Y(_05037_)
  );
  XNOR2X1 _12970_ (
    .A(_04961_),
    .B(_04962_),
    .Y(_05038_)
  );
  NAND2X1 _12971_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05038_),
    .Y(_05039_)
  );
  NAND2X1 _12972_ (
    .A(_05009_),
    .B(_05039_),
    .Y(_05040_)
  );
  OR2X1 _12973_ (
    .A(_05325_),
    .B(_05040_),
    .Y(_05041_)
  );
  XNOR2X1 _12974_ (
    .A(_05325_),
    .B(_05040_),
    .Y(_05042_)
  );
  NOR2X1 _12975_ (
    .A(_05334_),
    .B(_04637_),
    .Y(_05043_)
  );
  AOI21X1 _12976_ (
    .A(_05334_),
    .B(_05008_),
    .C(_05043_),
    .Y(_05044_)
  );
  AND2X1 _12977_ (
    .A( multiplier_0.reshi_7_ ),
    .B(_05044_),
    .Y(_05045_)
  );
  XOR2X1 _12978_ (
    .A( multiplier_0.reshi_7_ ),
    .B(_05044_),
    .Y(_05046_)
  );
  MUX2X1 _12979_ (
    .A(_05899_),
    .B(_04992_),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05047_)
  );
  NAND2X1 _12980_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_05047_),
    .Y(_05048_)
  );
  XNOR2X1 _12981_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_05047_),
    .Y(_05049_)
  );
  MUX2X1 _12982_ (
    .A(_05905_),
    .B(_05013_),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05050_)
  );
  NOR2X1 _12983_ (
    .A(_05326_),
    .B(_05050_),
    .Y(_05051_)
  );
  NAND2X1 _12984_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05911_),
    .Y(_05052_)
  );
  OAI21X1 _12985_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05018_),
    .C(_05052_),
    .Y(_05053_)
  );
  NOR2X1 _12986_ (
    .A(_05327_),
    .B(_05053_),
    .Y(_05054_)
  );
  OR2X1 _12987_ (
    .A(_05327_),
    .B(_05053_),
    .Y(_05055_)
  );
  AND2X1 _12988_ (
    .A(_05327_),
    .B(_05053_),
    .Y(_05056_)
  );
  NOR2X1 _12989_ (
    .A(_05054_),
    .B(_05056_),
    .Y(_05057_)
  );
  NAND2X1 _12990_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05916_),
    .Y(_05058_)
  );
  OAI21X1 _12991_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_05022_),
    .C(_05058_),
    .Y(_05059_)
  );
  NOR2X1 _12992_ (
    .A(_05328_),
    .B(_05059_),
    .Y(_05060_)
  );
  MUX2X1 _12993_ (
    .A(_05924_),
    .B(_05027_),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05061_)
  );
  NOR2X1 _12994_ (
    .A(_05329_),
    .B(_05061_),
    .Y(_05062_)
  );
  OR2X1 _12995_ (
    .A(_05329_),
    .B(_05061_),
    .Y(_05063_)
  );
  AND2X1 _12996_ (
    .A(_05329_),
    .B(_05061_),
    .Y(_05064_)
  );
  NOR2X1 _12997_ (
    .A(_05062_),
    .B(_05064_),
    .Y(_05065_)
  );
  MUX2X1 _12998_ (
    .A(_05931_),
    .B(_05032_),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05066_)
  );
  AND2X1 _12999_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_05066_),
    .Y(_05067_)
  );
  NAND2X1 _13000_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_05066_),
    .Y(_05068_)
  );
  MUX2X1 _13001_ (
    .A(_05939_),
    .B(_05038_),
    .S( multiplier_0.cycle_0_ ),
    .Y(_05069_)
  );
  NAND2X1 _13002_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_05069_),
    .Y(_05070_)
  );
  AOI21X1 _13003_ (
    .A(_05990_),
    .B(_04641_),
    .C(_04640_),
    .Y(_05071_)
  );
  XNOR2X1 _13004_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_05069_),
    .Y(_05072_)
  );
  OAI21X1 _13005_ (
    .A(_05071_),
    .B(_05072_),
    .C(_05070_),
    .Y(_05073_)
  );
  OR2X1 _13006_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_05066_),
    .Y(_05074_)
  );
  NAND2X1 _13007_ (
    .A(_05068_),
    .B(_05074_),
    .Y(_05075_)
  );
  AOI21X1 _13008_ (
    .A(_05073_),
    .B(_05074_),
    .C(_05067_),
    .Y(_05076_)
  );
  OAI21X1 _13009_ (
    .A(_05064_),
    .B(_05076_),
    .C(_05063_),
    .Y(_05077_)
  );
  XNOR2X1 _13010_ (
    .A( multiplier_0.reshi_3_ ),
    .B(_05059_),
    .Y(_05078_)
  );
  AOI21X1 _13011_ (
    .A(_05077_),
    .B(_05078_),
    .C(_05060_),
    .Y(_05079_)
  );
  OAI21X1 _13012_ (
    .A(_05056_),
    .B(_05079_),
    .C(_05055_),
    .Y(_05080_)
  );
  XNOR2X1 _13013_ (
    .A( multiplier_0.reshi_5_ ),
    .B(_05050_),
    .Y(_05081_)
  );
  AOI21X1 _13014_ (
    .A(_05080_),
    .B(_05081_),
    .C(_05051_),
    .Y(_05082_)
  );
  OAI21X1 _13015_ (
    .A(_05049_),
    .B(_05082_),
    .C(_05048_),
    .Y(_05083_)
  );
  AOI21X1 _13016_ (
    .A(_05046_),
    .B(_05083_),
    .C(_05045_),
    .Y(_05084_)
  );
  OAI21X1 _13017_ (
    .A(_05042_),
    .B(_05084_),
    .C(_05041_),
    .Y(_05085_)
  );
  OAI21X1 _13018_ (
    .A(_05036_),
    .B(_05085_),
    .C(_05037_),
    .Y(_05086_)
  );
  OAI21X1 _13019_ (
    .A(_05031_),
    .B(_05086_),
    .C(_05030_),
    .Y(_05087_)
  );
  AOI21X1 _13020_ (
    .A(_05024_),
    .B(_05087_),
    .C(_05026_),
    .Y(_05088_)
  );
  OAI21X1 _13021_ (
    .A(_05021_),
    .B(_05088_),
    .C(_05020_),
    .Y(_05089_)
  );
  AOI21X1 _13022_ (
    .A(_05015_),
    .B(_05089_),
    .C(_05017_),
    .Y(_05090_)
  );
  OAI21X1 _13023_ (
    .A(_05012_),
    .B(_05090_),
    .C(_05011_),
    .Y(_05091_)
  );
  AOI21X1 _13024_ (
    .A(_05332_),
    .B(_05334_),
    .C(_05008_),
    .Y(_05092_)
  );
  XNOR2X1 _13025_ (
    .A( multiplier_0.reshi_15_ ),
    .B(_05092_),
    .Y(_05093_)
  );
  INVX1 _13026_ (
    .A(_05093_),
    .Y(_05094_)
  );
  NAND2X1 _13027_ (
    .A(_05091_),
    .B(_05094_),
    .Y(_05095_)
  );
  XNOR2X1 _13028_ (
    .A(_05091_),
    .B(_05094_),
    .Y(_05096_)
  );
  AOI21X1 _13029_ (
    .A(_05361_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05097_)
  );
  OAI21X1 _13030_ (
    .A(_04716_),
    .B(_05096_),
    .C(_05097_),
    .Y(_05098_)
  );
  OAI21X1 _13031_ (
    .A( multiplier_0.reshi_15_ ),
    .B(_04718_),
    .C(_05098_),
    .Y(_05099_)
  );
  INVX1 _13032_ (
    .A(_05099_),
    .Y(_04553_)
  );
  XNOR2X1 _13033_ (
    .A(_05012_),
    .B(_05090_),
    .Y(_05100_)
  );
  AOI21X1 _13034_ (
    .A(_05364_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05101_)
  );
  OAI21X1 _13035_ (
    .A(_04716_),
    .B(_05100_),
    .C(_05101_),
    .Y(_05102_)
  );
  OAI21X1 _13036_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_04718_),
    .C(_05102_),
    .Y(_05103_)
  );
  INVX1 _13037_ (
    .A(_05103_),
    .Y(_04552_)
  );
  NAND2X1 _13038_ (
    .A(_05015_),
    .B(_05016_),
    .Y(_05104_)
  );
  XOR2X1 _13039_ (
    .A(_05089_),
    .B(_05104_),
    .Y(_05105_)
  );
  AOI21X1 _13040_ (
    .A(_05367_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05106_)
  );
  OAI21X1 _13041_ (
    .A(_04716_),
    .B(_05105_),
    .C(_05106_),
    .Y(_05107_)
  );
  OAI21X1 _13042_ (
    .A( multiplier_0.reshi_13_ ),
    .B(_04718_),
    .C(_05107_),
    .Y(_05108_)
  );
  INVX1 _13043_ (
    .A(_05108_),
    .Y(_04551_)
  );
  XNOR2X1 _13044_ (
    .A(_05021_),
    .B(_05088_),
    .Y(_05109_)
  );
  AOI21X1 _13045_ (
    .A(_05370_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05110_)
  );
  OAI21X1 _13046_ (
    .A(_04716_),
    .B(_05109_),
    .C(_05110_),
    .Y(_05111_)
  );
  OAI21X1 _13047_ (
    .A( multiplier_0.reshi_12_ ),
    .B(_04718_),
    .C(_05111_),
    .Y(_05112_)
  );
  INVX1 _13048_ (
    .A(_05112_),
    .Y(_04550_)
  );
  NAND2X1 _13049_ (
    .A(_05024_),
    .B(_05025_),
    .Y(_05113_)
  );
  XOR2X1 _13050_ (
    .A(_05087_),
    .B(_05113_),
    .Y(_05114_)
  );
  AOI21X1 _13051_ (
    .A(_05373_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05115_)
  );
  OAI21X1 _13052_ (
    .A(_04716_),
    .B(_05114_),
    .C(_05115_),
    .Y(_05116_)
  );
  OAI21X1 _13053_ (
    .A( multiplier_0.reshi_11_ ),
    .B(_04718_),
    .C(_05116_),
    .Y(_05117_)
  );
  INVX1 _13054_ (
    .A(_05117_),
    .Y(_04549_)
  );
  XNOR2X1 _13055_ (
    .A(_05031_),
    .B(_05086_),
    .Y(_05118_)
  );
  AOI21X1 _13056_ (
    .A(_05376_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05119_)
  );
  OAI21X1 _13057_ (
    .A(_04716_),
    .B(_05118_),
    .C(_05119_),
    .Y(_05120_)
  );
  OAI21X1 _13058_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_04718_),
    .C(_05120_),
    .Y(_05121_)
  );
  INVX1 _13059_ (
    .A(_05121_),
    .Y(_04548_)
  );
  NAND2X1 _13060_ (
    .A(_05035_),
    .B(_05037_),
    .Y(_05122_)
  );
  XOR2X1 _13061_ (
    .A(_05085_),
    .B(_05122_),
    .Y(_05123_)
  );
  AOI21X1 _13062_ (
    .A(_05379_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05124_)
  );
  OAI21X1 _13063_ (
    .A(_04716_),
    .B(_05123_),
    .C(_05124_),
    .Y(_05125_)
  );
  OAI21X1 _13064_ (
    .A( multiplier_0.reshi_9_ ),
    .B(_04718_),
    .C(_05125_),
    .Y(_05126_)
  );
  INVX1 _13065_ (
    .A(_05126_),
    .Y(_04547_)
  );
  XNOR2X1 _13066_ (
    .A(_05042_),
    .B(_05084_),
    .Y(_05127_)
  );
  AOI21X1 _13067_ (
    .A(_05382_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05128_)
  );
  OAI21X1 _13068_ (
    .A(_04716_),
    .B(_05127_),
    .C(_05128_),
    .Y(_05129_)
  );
  OAI21X1 _13069_ (
    .A( multiplier_0.reshi_8_ ),
    .B(_04718_),
    .C(_05129_),
    .Y(_05130_)
  );
  INVX1 _13070_ (
    .A(_05130_),
    .Y(_04546_)
  );
  XNOR2X1 _13071_ (
    .A(_05046_),
    .B(_05083_),
    .Y(_05131_)
  );
  AOI21X1 _13072_ (
    .A(_06288_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05132_)
  );
  OAI21X1 _13073_ (
    .A(_04716_),
    .B(_05131_),
    .C(_05132_),
    .Y(_05133_)
  );
  OAI21X1 _13074_ (
    .A( multiplier_0.reshi_7_ ),
    .B(_04718_),
    .C(_05133_),
    .Y(_05134_)
  );
  INVX1 _13075_ (
    .A(_05134_),
    .Y(_04545_)
  );
  XNOR2X1 _13076_ (
    .A(_05049_),
    .B(_05082_),
    .Y(_05135_)
  );
  AOI21X1 _13077_ (
    .A(_06287_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05136_)
  );
  OAI21X1 _13078_ (
    .A(_04716_),
    .B(_05135_),
    .C(_05136_),
    .Y(_05137_)
  );
  OAI21X1 _13079_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_04718_),
    .C(_05137_),
    .Y(_05138_)
  );
  INVX1 _13080_ (
    .A(_05138_),
    .Y(_04544_)
  );
  XNOR2X1 _13081_ (
    .A(_05080_),
    .B(_05081_),
    .Y(_05139_)
  );
  AOI21X1 _13082_ (
    .A(_06286_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05140_)
  );
  OAI21X1 _13083_ (
    .A(_04716_),
    .B(_05139_),
    .C(_05140_),
    .Y(_05141_)
  );
  OAI21X1 _13084_ (
    .A( multiplier_0.reshi_5_ ),
    .B(_04718_),
    .C(_05141_),
    .Y(_05142_)
  );
  INVX1 _13085_ (
    .A(_05142_),
    .Y(_04543_)
  );
  XOR2X1 _13086_ (
    .A(_05057_),
    .B(_05079_),
    .Y(_05143_)
  );
  AOI21X1 _13087_ (
    .A(_06285_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05144_)
  );
  OAI21X1 _13088_ (
    .A(_04716_),
    .B(_05143_),
    .C(_05144_),
    .Y(_05145_)
  );
  OAI21X1 _13089_ (
    .A( multiplier_0.reshi_4_ ),
    .B(_04718_),
    .C(_05145_),
    .Y(_05146_)
  );
  INVX1 _13090_ (
    .A(_05146_),
    .Y(_04542_)
  );
  XNOR2X1 _13091_ (
    .A(_05077_),
    .B(_05078_),
    .Y(_05147_)
  );
  AOI21X1 _13092_ (
    .A(_06284_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05148_)
  );
  OAI21X1 _13093_ (
    .A(_04716_),
    .B(_05147_),
    .C(_05148_),
    .Y(_05149_)
  );
  OAI21X1 _13094_ (
    .A( multiplier_0.reshi_3_ ),
    .B(_04718_),
    .C(_05149_),
    .Y(_05150_)
  );
  INVX1 _13095_ (
    .A(_05150_),
    .Y(_04541_)
  );
  XOR2X1 _13096_ (
    .A(_05065_),
    .B(_05076_),
    .Y(_05151_)
  );
  AOI21X1 _13097_ (
    .A(_06283_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05152_)
  );
  OAI21X1 _13098_ (
    .A(_04716_),
    .B(_05151_),
    .C(_05152_),
    .Y(_05153_)
  );
  OAI21X1 _13099_ (
    .A( multiplier_0.reshi_2_ ),
    .B(_04718_),
    .C(_05153_),
    .Y(_05154_)
  );
  INVX1 _13100_ (
    .A(_05154_),
    .Y(_04540_)
  );
  XOR2X1 _13101_ (
    .A(_05073_),
    .B(_05075_),
    .Y(_05155_)
  );
  AOI21X1 _13102_ (
    .A(_06282_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05156_)
  );
  OAI21X1 _13103_ (
    .A(_04716_),
    .B(_05155_),
    .C(_05156_),
    .Y(_05157_)
  );
  OAI21X1 _13104_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_04718_),
    .C(_05157_),
    .Y(_05158_)
  );
  INVX1 _13105_ (
    .A(_05158_),
    .Y(_04539_)
  );
  XNOR2X1 _13106_ (
    .A(_05071_),
    .B(_05072_),
    .Y(_05159_)
  );
  AOI21X1 _13107_ (
    .A(_06275_),
    .B(_04715_),
    .C(_04717_),
    .Y(_05160_)
  );
  OAI21X1 _13108_ (
    .A(_04716_),
    .B(_05159_),
    .C(_05160_),
    .Y(_05161_)
  );
  OAI21X1 _13109_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_04718_),
    .C(_05161_),
    .Y(_05162_)
  );
  INVX1 _13110_ (
    .A(_05162_),
    .Y(_04538_)
  );
  OAI21X1 _13111_ (
    .A(_05351_),
    .B(_05393_),
    .C(_05411_),
    .Y(_05163_)
  );
  NOR2X1 _13112_ (
    .A(_05332_),
    .B(_05096_),
    .Y(_05164_)
  );
  NOR2X1 _13113_ (
    .A( multiplier_0.op2_wr ),
    .B(_05411_),
    .Y(_05165_)
  );
  NAND2X1 _13114_ (
    .A(_05164_),
    .B(_05165_),
    .Y(_05166_)
  );
  OAI21X1 _13115_ (
    .A(_05330_),
    .B(_05163_),
    .C(_05166_),
    .Y(_04537_)
  );
  AOI21X1 _13116_ (
    .A( multiplier_0.reshi_15_ ),
    .B(_05092_),
    .C( multiplier_0.sumext_0_ ),
    .Y(_05167_)
  );
  AOI21X1 _13117_ (
    .A(_05095_),
    .B(_05167_),
    .C( multiplier_0.sign_sel ),
    .Y(_05168_)
  );
  OAI21X1 _13118_ (
    .A(_05164_),
    .B(_05168_),
    .C(_05165_),
    .Y(_05169_)
  );
  OAI21X1 _13119_ (
    .A(_05331_),
    .B(_05163_),
    .C(_05169_),
    .Y(_04536_)
  );
  MUX2X1 _13120_ (
    .A( multiplier_0.sign_sel ),
    .B(_06262_),
    .S(_05359_),
    .Y(_05170_)
  );
  INVX1 _13121_ (
    .A(_05170_),
    .Y(_04535_)
  );
  MUX2X1 _13122_ (
    .A( multiplier_0.acc_sel ),
    .B(_06266_),
    .S(_05359_),
    .Y(_05171_)
  );
  INVX1 _13123_ (
    .A(_05171_),
    .Y(_04534_)
  );
  OAI21X1 _13124_ (
    .A(_05332_),
    .B(_05096_),
    .C( multiplier_0.cycle_1_ ),
    .Y(_05172_)
  );
  NOR2X1 _13125_ (
    .A(_05168_),
    .B(_05172_),
    .Y(_05173_)
  );
  NAND2X1 _13126_ (
    .A(_05340_),
    .B(_05350_),
    .Y(_05174_)
  );
  NAND3X1 _13127_ (
    .A(_06262_),
    .B(_05340_),
    .C(_05350_),
    .Y(_05175_)
  );
  NOR2X1 _13128_ (
    .A(_04713_),
    .B(_05175_),
    .Y(_05176_)
  );
  OAI21X1 _13129_ (
    .A( multiplier_0.sumext_0_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05176_),
    .Y(_05177_)
  );
  NOR2X1 _13130_ (
    .A(_04714_),
    .B(_05174_),
    .Y(_05178_)
  );
  OAI21X1 _13131_ (
    .A( multiplier_0.reshi_0_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05179_)
  );
  AOI21X1 _13132_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05159_),
    .C(_05179_),
    .Y(_05180_)
  );
  NOR2X1 _13133_ (
    .A(_05392_),
    .B(_05175_),
    .Y(_05181_)
  );
  INVX1 _13134_ (
    .A(_05181_),
    .Y(_05182_)
  );
  NAND2X1 _13135_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04709_),
    .Y(_05183_)
  );
  OAI21X1 _13136_ (
    .A( multiplier_0.reslo_0_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05183_),
    .Y(_05184_)
  );
  NOR2X1 _13137_ (
    .A(_05393_),
    .B(_05174_),
    .Y(_05185_)
  );
  NOR2X1 _13138_ (
    .A(_06267_),
    .B(_05174_),
    .Y(_05186_)
  );
  AOI22X1 _13139_ (
    .A( multiplier_0.op2_0_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_0_ ),
    .Y(_05187_)
  );
  OAI21X1 _13140_ (
    .A(_05182_),
    .B(_05184_),
    .C(_05187_),
    .Y(_05188_)
  );
  NOR2X1 _13141_ (
    .A(_05180_),
    .B(_05188_),
    .Y(_05189_)
  );
  OAI21X1 _13142_ (
    .A(_05173_),
    .B(_05177_),
    .C(_05189_),
    .Y( multiplier_0.per_dout_0_ )
  );
  OAI21X1 _13143_ (
    .A( multiplier_0.sumext_10_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05176_),
    .Y(_05190_)
  );
  INVX1 _13144_ (
    .A(_05190_),
    .Y(_05191_)
  );
  OAI21X1 _13145_ (
    .A(_05333_),
    .B(_05164_),
    .C(_05191_),
    .Y(_05192_)
  );
  OAI21X1 _13146_ (
    .A( multiplier_0.reshi_1_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05193_)
  );
  AOI21X1 _13147_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05155_),
    .C(_05193_),
    .Y(_05194_)
  );
  AND2X1 _13148_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04704_),
    .Y(_05195_)
  );
  OAI21X1 _13149_ (
    .A( multiplier_0.reslo_1_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05196_)
  );
  AOI22X1 _13150_ (
    .A( multiplier_0.op2_1_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_1_ ),
    .Y(_05197_)
  );
  OAI21X1 _13151_ (
    .A(_05195_),
    .B(_05196_),
    .C(_05197_),
    .Y(_05198_)
  );
  NOR2X1 _13152_ (
    .A(_05194_),
    .B(_05198_),
    .Y(_05199_)
  );
  NAND2X1 _13153_ (
    .A(_05192_),
    .B(_05199_),
    .Y( multiplier_0.per_dout_1_ )
  );
  OAI21X1 _13154_ (
    .A( multiplier_0.reshi_2_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05200_)
  );
  AOI21X1 _13155_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05151_),
    .C(_05200_),
    .Y(_05201_)
  );
  AND2X1 _13156_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04700_),
    .Y(_05202_)
  );
  OAI21X1 _13157_ (
    .A( multiplier_0.reslo_2_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05203_)
  );
  AOI22X1 _13158_ (
    .A( multiplier_0.op2_2_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_2_ ),
    .Y(_05204_)
  );
  OAI21X1 _13159_ (
    .A(_05202_),
    .B(_05203_),
    .C(_05204_),
    .Y(_05205_)
  );
  NOR2X1 _13160_ (
    .A(_05201_),
    .B(_05205_),
    .Y(_05206_)
  );
  NAND2X1 _13161_ (
    .A(_05192_),
    .B(_05206_),
    .Y( multiplier_0.per_dout_2_ )
  );
  OAI21X1 _13162_ (
    .A( multiplier_0.reshi_3_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05207_)
  );
  AOI21X1 _13163_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05147_),
    .C(_05207_),
    .Y(_05208_)
  );
  NOR2X1 _13164_ (
    .A(_05333_),
    .B(_04695_),
    .Y(_05209_)
  );
  OAI21X1 _13165_ (
    .A( multiplier_0.reslo_3_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05210_)
  );
  AOI22X1 _13166_ (
    .A( multiplier_0.op2_3_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_3_ ),
    .Y(_05211_)
  );
  OAI21X1 _13167_ (
    .A(_05209_),
    .B(_05210_),
    .C(_05211_),
    .Y(_05212_)
  );
  NOR2X1 _13168_ (
    .A(_05208_),
    .B(_05212_),
    .Y(_05213_)
  );
  NAND2X1 _13169_ (
    .A(_05192_),
    .B(_05213_),
    .Y( multiplier_0.per_dout_3_ )
  );
  OAI21X1 _13170_ (
    .A( multiplier_0.reshi_4_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05214_)
  );
  AOI21X1 _13171_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05143_),
    .C(_05214_),
    .Y(_05215_)
  );
  NOR2X1 _13172_ (
    .A(_05333_),
    .B(_04690_),
    .Y(_05216_)
  );
  OAI21X1 _13173_ (
    .A( multiplier_0.reslo_4_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05217_)
  );
  AOI22X1 _13174_ (
    .A( multiplier_0.op2_4_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_4_ ),
    .Y(_05218_)
  );
  OAI21X1 _13175_ (
    .A(_05216_),
    .B(_05217_),
    .C(_05218_),
    .Y(_05219_)
  );
  NOR2X1 _13176_ (
    .A(_05215_),
    .B(_05219_),
    .Y(_05220_)
  );
  NAND2X1 _13177_ (
    .A(_05192_),
    .B(_05220_),
    .Y( multiplier_0.per_dout_4_ )
  );
  OAI21X1 _13178_ (
    .A( multiplier_0.reshi_5_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05221_)
  );
  AOI21X1 _13179_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05139_),
    .C(_05221_),
    .Y(_05222_)
  );
  NOR2X1 _13180_ (
    .A(_05333_),
    .B(_04685_),
    .Y(_05223_)
  );
  OAI21X1 _13181_ (
    .A( multiplier_0.reslo_5_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05224_)
  );
  AOI22X1 _13182_ (
    .A( multiplier_0.op2_5_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_5_ ),
    .Y(_05225_)
  );
  OAI21X1 _13183_ (
    .A(_05223_),
    .B(_05224_),
    .C(_05225_),
    .Y(_05226_)
  );
  NOR2X1 _13184_ (
    .A(_05222_),
    .B(_05226_),
    .Y(_05227_)
  );
  NAND2X1 _13185_ (
    .A(_05192_),
    .B(_05227_),
    .Y( multiplier_0.per_dout_5_ )
  );
  OAI21X1 _13186_ (
    .A( multiplier_0.reshi_6_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05228_)
  );
  AOI21X1 _13187_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05135_),
    .C(_05228_),
    .Y(_05229_)
  );
  AND2X1 _13188_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04681_),
    .Y(_05230_)
  );
  OAI21X1 _13189_ (
    .A( multiplier_0.reslo_6_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05231_)
  );
  AOI22X1 _13190_ (
    .A( multiplier_0.op2_6_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_6_ ),
    .Y(_05232_)
  );
  OAI21X1 _13191_ (
    .A(_05230_),
    .B(_05231_),
    .C(_05232_),
    .Y(_05233_)
  );
  NOR2X1 _13192_ (
    .A(_05229_),
    .B(_05233_),
    .Y(_05234_)
  );
  NAND2X1 _13193_ (
    .A(_05192_),
    .B(_05234_),
    .Y( multiplier_0.per_dout_6_ )
  );
  OAI21X1 _13194_ (
    .A( multiplier_0.reshi_7_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05235_)
  );
  AOI21X1 _13195_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05131_),
    .C(_05235_),
    .Y(_05236_)
  );
  NOR2X1 _13196_ (
    .A(_05333_),
    .B(_04676_),
    .Y(_05237_)
  );
  OAI21X1 _13197_ (
    .A( multiplier_0.reslo_7_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05238_)
  );
  AOI22X1 _13198_ (
    .A( multiplier_0.op2_7_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_7_ ),
    .Y(_05239_)
  );
  OAI21X1 _13199_ (
    .A(_05237_),
    .B(_05238_),
    .C(_05239_),
    .Y(_05240_)
  );
  NOR2X1 _13200_ (
    .A(_05236_),
    .B(_05240_),
    .Y(_05241_)
  );
  NAND2X1 _13201_ (
    .A(_05192_),
    .B(_05241_),
    .Y( multiplier_0.per_dout_7_ )
  );
  OAI21X1 _13202_ (
    .A( multiplier_0.reshi_8_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05242_)
  );
  AOI21X1 _13203_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05127_),
    .C(_05242_),
    .Y(_05243_)
  );
  AND2X1 _13204_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04672_),
    .Y(_05244_)
  );
  OAI21X1 _13205_ (
    .A( multiplier_0.reslo_8_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05245_)
  );
  AOI22X1 _13206_ (
    .A( multiplier_0.op2_8_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_8_ ),
    .Y(_05246_)
  );
  OAI21X1 _13207_ (
    .A(_05244_),
    .B(_05245_),
    .C(_05246_),
    .Y(_05247_)
  );
  NOR2X1 _13208_ (
    .A(_05243_),
    .B(_05247_),
    .Y(_05248_)
  );
  NAND2X1 _13209_ (
    .A(_05192_),
    .B(_05248_),
    .Y( multiplier_0.per_dout_8_ )
  );
  OAI21X1 _13210_ (
    .A( multiplier_0.reshi_9_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05249_)
  );
  AOI21X1 _13211_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05123_),
    .C(_05249_),
    .Y(_05250_)
  );
  AND2X1 _13212_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04668_),
    .Y(_05251_)
  );
  OAI21X1 _13213_ (
    .A( multiplier_0.reslo_9_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05252_)
  );
  AOI22X1 _13214_ (
    .A( multiplier_0.op2_9_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_9_ ),
    .Y(_05253_)
  );
  OAI21X1 _13215_ (
    .A(_05251_),
    .B(_05252_),
    .C(_05253_),
    .Y(_05254_)
  );
  NOR2X1 _13216_ (
    .A(_05250_),
    .B(_05254_),
    .Y(_05255_)
  );
  NAND2X1 _13217_ (
    .A(_05192_),
    .B(_05255_),
    .Y( multiplier_0.per_dout_9_ )
  );
  OAI21X1 _13218_ (
    .A( multiplier_0.reshi_10_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05256_)
  );
  AOI21X1 _13219_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05118_),
    .C(_05256_),
    .Y(_05257_)
  );
  AND2X1 _13220_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04664_),
    .Y(_05258_)
  );
  OAI21X1 _13221_ (
    .A( multiplier_0.reslo_10_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05259_)
  );
  AOI22X1 _13222_ (
    .A( multiplier_0.op2_10_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_10_ ),
    .Y(_05260_)
  );
  OAI21X1 _13223_ (
    .A(_05258_),
    .B(_05259_),
    .C(_05260_),
    .Y(_05261_)
  );
  NOR2X1 _13224_ (
    .A(_05257_),
    .B(_05261_),
    .Y(_05262_)
  );
  NAND2X1 _13225_ (
    .A(_05192_),
    .B(_05262_),
    .Y( multiplier_0.per_dout_10_ )
  );
  OAI21X1 _13226_ (
    .A( multiplier_0.reshi_11_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05263_)
  );
  AOI21X1 _13227_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05114_),
    .C(_05263_),
    .Y(_05264_)
  );
  AND2X1 _13228_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04660_),
    .Y(_05265_)
  );
  OAI21X1 _13229_ (
    .A( multiplier_0.reslo_11_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05266_)
  );
  AOI22X1 _13230_ (
    .A( multiplier_0.op2_11_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_11_ ),
    .Y(_05267_)
  );
  OAI21X1 _13231_ (
    .A(_05265_),
    .B(_05266_),
    .C(_05267_),
    .Y(_05268_)
  );
  NOR2X1 _13232_ (
    .A(_05264_),
    .B(_05268_),
    .Y(_05269_)
  );
  NAND2X1 _13233_ (
    .A(_05192_),
    .B(_05269_),
    .Y( multiplier_0.per_dout_11_ )
  );
  OAI21X1 _13234_ (
    .A( multiplier_0.reshi_12_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05270_)
  );
  AOI21X1 _13235_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05109_),
    .C(_05270_),
    .Y(_05271_)
  );
  AND2X1 _13236_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04656_),
    .Y(_05272_)
  );
  OAI21X1 _13237_ (
    .A( multiplier_0.reslo_12_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05273_)
  );
  AOI22X1 _13238_ (
    .A( multiplier_0.op2_12_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_12_ ),
    .Y(_05274_)
  );
  OAI21X1 _13239_ (
    .A(_05272_),
    .B(_05273_),
    .C(_05274_),
    .Y(_05275_)
  );
  NOR2X1 _13240_ (
    .A(_05271_),
    .B(_05275_),
    .Y(_05276_)
  );
  NAND2X1 _13241_ (
    .A(_05192_),
    .B(_05276_),
    .Y( multiplier_0.per_dout_12_ )
  );
  OAI21X1 _13242_ (
    .A( multiplier_0.reshi_13_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05277_)
  );
  AOI21X1 _13243_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05105_),
    .C(_05277_),
    .Y(_05278_)
  );
  AND2X1 _13244_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04652_),
    .Y(_05279_)
  );
  OAI21X1 _13245_ (
    .A( multiplier_0.reslo_13_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05280_)
  );
  AOI22X1 _13246_ (
    .A( multiplier_0.op2_13_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_13_ ),
    .Y(_05281_)
  );
  OAI21X1 _13247_ (
    .A(_05279_),
    .B(_05280_),
    .C(_05281_),
    .Y(_05282_)
  );
  NOR2X1 _13248_ (
    .A(_05278_),
    .B(_05282_),
    .Y(_05283_)
  );
  NAND2X1 _13249_ (
    .A(_05192_),
    .B(_05283_),
    .Y( multiplier_0.per_dout_13_ )
  );
  OAI21X1 _13250_ (
    .A( multiplier_0.reshi_14_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05284_)
  );
  AOI21X1 _13251_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05100_),
    .C(_05284_),
    .Y(_05285_)
  );
  AOI21X1 _13252_ (
    .A(_05989_),
    .B(_04647_),
    .C(_05333_),
    .Y(_05286_)
  );
  OAI21X1 _13253_ (
    .A( multiplier_0.reslo_14_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05287_)
  );
  AOI22X1 _13254_ (
    .A( multiplier_0.op2_14_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_14_ ),
    .Y(_05288_)
  );
  OAI21X1 _13255_ (
    .A(_05286_),
    .B(_05287_),
    .C(_05288_),
    .Y(_05289_)
  );
  NOR2X1 _13256_ (
    .A(_05285_),
    .B(_05289_),
    .Y(_05290_)
  );
  NAND2X1 _13257_ (
    .A(_05192_),
    .B(_05290_),
    .Y( multiplier_0.per_dout_14_ )
  );
  OAI21X1 _13258_ (
    .A( multiplier_0.reshi_15_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05178_),
    .Y(_05291_)
  );
  AOI21X1 _13259_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_05096_),
    .C(_05291_),
    .Y(_05292_)
  );
  AND2X1 _13260_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04643_),
    .Y(_05293_)
  );
  OAI21X1 _13261_ (
    .A( multiplier_0.reslo_15_ ),
    .B( multiplier_0.cycle_1_ ),
    .C(_05181_),
    .Y(_05294_)
  );
  AOI22X1 _13262_ (
    .A( multiplier_0.op2_15_ ),
    .B(_05185_),
    .C(_05186_),
    .D( multiplier_0.op1_15_ ),
    .Y(_05295_)
  );
  OAI21X1 _13263_ (
    .A(_05293_),
    .B(_05294_),
    .C(_05295_),
    .Y(_05296_)
  );
  NOR2X1 _13264_ (
    .A(_05292_),
    .B(_05296_),
    .Y(_05297_)
  );
  NAND2X1 _13265_ (
    .A(_05192_),
    .B(_05297_),
    .Y( multiplier_0.per_dout_15_ )
  );
  INVX1 _13266_ (
    .A(_06327_),
    .Y(_04465_)
  );
  INVX1 _13267_ (
    .A(_06327_),
    .Y(_04466_)
  );
  INVX1 _13268_ (
    .A(_06327_),
    .Y(_04467_)
  );
  INVX1 _13269_ (
    .A(_06327_),
    .Y(_04468_)
  );
  INVX1 _13270_ (
    .A(_06327_),
    .Y(_04469_)
  );
  INVX1 _13271_ (
    .A(_06327_),
    .Y(_04470_)
  );
  INVX1 _13272_ (
    .A(_06327_),
    .Y(_04471_)
  );
  INVX1 _13273_ (
    .A(_06327_),
    .Y(_04472_)
  );
  INVX1 _13274_ (
    .A(_06327_),
    .Y(_04473_)
  );
  INVX1 _13275_ (
    .A(_06327_),
    .Y(_04474_)
  );
  INVX1 _13276_ (
    .A(_06327_),
    .Y(_04475_)
  );
  INVX1 _13277_ (
    .A(_06327_),
    .Y(_04476_)
  );
  INVX1 _13278_ (
    .A(_06327_),
    .Y(_04477_)
  );
  INVX1 _13279_ (
    .A(_06327_),
    .Y(_04478_)
  );
  INVX1 _13280_ (
    .A(_06327_),
    .Y(_04479_)
  );
  INVX1 _13281_ (
    .A(_06327_),
    .Y(_04480_)
  );
  INVX1 _13282_ (
    .A(_06327_),
    .Y(_04481_)
  );
  INVX1 _13283_ (
    .A(_06327_),
    .Y(_04482_)
  );
  INVX1 _13284_ (
    .A(_06327_),
    .Y(_04483_)
  );
  INVX1 _13285_ (
    .A(_06327_),
    .Y(_04484_)
  );
  INVX1 _13286_ (
    .A(_06327_),
    .Y(_04485_)
  );
  INVX1 _13287_ (
    .A(_06327_),
    .Y(_04486_)
  );
  INVX1 _13288_ (
    .A(_06327_),
    .Y(_04487_)
  );
  INVX1 _13289_ (
    .A(_06327_),
    .Y(_04488_)
  );
  INVX1 _13290_ (
    .A(_06327_),
    .Y(_04489_)
  );
  INVX1 _13291_ (
    .A(_06327_),
    .Y(_04490_)
  );
  INVX1 _13292_ (
    .A(_06327_),
    .Y(_04491_)
  );
  INVX1 _13293_ (
    .A(_06327_),
    .Y(_04492_)
  );
  INVX1 _13294_ (
    .A(_06327_),
    .Y(_04493_)
  );
  INVX1 _13295_ (
    .A(_06327_),
    .Y(_04494_)
  );
  INVX1 _13296_ (
    .A(_06327_),
    .Y(_04495_)
  );
  INVX1 _13297_ (
    .A(_06327_),
    .Y(_04496_)
  );
  INVX1 _13298_ (
    .A(_06327_),
    .Y(_04497_)
  );
  INVX1 _13299_ (
    .A(_06327_),
    .Y(_04498_)
  );
  INVX1 _13300_ (
    .A(_06327_),
    .Y(_04499_)
  );
  INVX1 _13301_ (
    .A(_06327_),
    .Y(_04500_)
  );
  INVX1 _13302_ (
    .A(_06327_),
    .Y(_04501_)
  );
  INVX1 _13303_ (
    .A(_06327_),
    .Y(_04502_)
  );
  INVX1 _13304_ (
    .A(_06327_),
    .Y(_04503_)
  );
  INVX1 _13305_ (
    .A(_06327_),
    .Y(_04504_)
  );
  INVX1 _13306_ (
    .A(_06327_),
    .Y(_04505_)
  );
  INVX1 _13307_ (
    .A(_06327_),
    .Y(_04506_)
  );
  INVX1 _13308_ (
    .A(_06327_),
    .Y(_04507_)
  );
  INVX1 _13309_ (
    .A(_06327_),
    .Y(_04508_)
  );
  INVX1 _13310_ (
    .A(_06327_),
    .Y(_04509_)
  );
  INVX1 _13311_ (
    .A(_06327_),
    .Y(_04510_)
  );
  INVX1 _13312_ (
    .A(_06327_),
    .Y(_04511_)
  );
  INVX1 _13313_ (
    .A(_06327_),
    .Y(_04512_)
  );
  INVX1 _13314_ (
    .A(_06327_),
    .Y(_04513_)
  );
  INVX1 _13315_ (
    .A(_06327_),
    .Y(_04514_)
  );
  INVX1 _13316_ (
    .A(_06327_),
    .Y(_04515_)
  );
  INVX1 _13317_ (
    .A(_06327_),
    .Y(_04516_)
  );
  INVX1 _13318_ (
    .A(_06327_),
    .Y(_04517_)
  );
  INVX1 _13319_ (
    .A(_06327_),
    .Y(_04518_)
  );
  INVX1 _13320_ (
    .A(_06327_),
    .Y(_04519_)
  );
  INVX1 _13321_ (
    .A(_06327_),
    .Y(_04520_)
  );
  INVX1 _13322_ (
    .A(_06327_),
    .Y(_04521_)
  );
  INVX1 _13323_ (
    .A(_06327_),
    .Y(_04522_)
  );
  INVX1 _13324_ (
    .A(_06327_),
    .Y(_04523_)
  );
  INVX1 _13325_ (
    .A(_06327_),
    .Y(_04524_)
  );
  INVX1 _13326_ (
    .A(_06327_),
    .Y(_04525_)
  );
  INVX1 _13327_ (
    .A(_06327_),
    .Y(_04526_)
  );
  INVX1 _13328_ (
    .A(_06327_),
    .Y(_04527_)
  );
  INVX1 _13329_ (
    .A(_06327_),
    .Y(_04528_)
  );
  INVX1 _13330_ (
    .A(_06327_),
    .Y(_04529_)
  );
  INVX1 _13331_ (
    .A(_06327_),
    .Y(_04530_)
  );
  INVX1 _13332_ (
    .A(_06327_),
    .Y(_04531_)
  );
  INVX1 _13333_ (
    .A(_06327_),
    .Y(_04532_)
  );
  INVX1 _13334_ (
    .A(_06327_),
    .Y(_04533_)
  );
  DFFSR _13335_ (
    .CLK(dco_clk),
    .D( multiplier_0.op2_wr ),
    .Q( multiplier_0.cycle_0_ ),
    .R(_04464_),
    .S(1'h1)
  );
  DFFSR _13336_ (
    .CLK(dco_clk),
    .D( multiplier_0.cycle_0_ ),
    .Q( multiplier_0.cycle_1_ ),
    .R(_04465_),
    .S(1'h1)
  );
  DFFSR _13337_ (
    .CLK(dco_clk),
    .D(_04534_),
    .Q( multiplier_0.acc_sel ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13338_ (
    .CLK(dco_clk),
    .D(_04535_),
    .Q( multiplier_0.sign_sel ),
    .R(_04467_),
    .S(1'h1)
  );
  DFFSR _13339_ (
    .CLK(dco_clk),
    .D(_04536_),
    .Q( multiplier_0.sumext_0_ ),
    .R(_04468_),
    .S(1'h1)
  );
  DFFSR _13340_ (
    .CLK(dco_clk),
    .D(_04537_),
    .Q( multiplier_0.sumext_10_ ),
    .R(_04469_),
    .S(1'h1)
  );
  DFFSR _13341_ (
    .CLK(dco_clk),
    .D(_04538_),
    .Q( multiplier_0.reshi_0_ ),
    .R(_04470_),
    .S(1'h1)
  );
  DFFSR _13342_ (
    .CLK(dco_clk),
    .D(_04539_),
    .Q( multiplier_0.reshi_1_ ),
    .R(_04471_),
    .S(1'h1)
  );
  DFFSR _13343_ (
    .CLK(dco_clk),
    .D(_04540_),
    .Q( multiplier_0.reshi_2_ ),
    .R(_04472_),
    .S(1'h1)
  );
  DFFSR _13344_ (
    .CLK(dco_clk),
    .D(_04541_),
    .Q( multiplier_0.reshi_3_ ),
    .R(_04473_),
    .S(1'h1)
  );
  DFFSR _13345_ (
    .CLK(dco_clk),
    .D(_04542_),
    .Q( multiplier_0.reshi_4_ ),
    .R(_04474_),
    .S(1'h1)
  );
  DFFSR _13346_ (
    .CLK(dco_clk),
    .D(_04543_),
    .Q( multiplier_0.reshi_5_ ),
    .R(_04475_),
    .S(1'h1)
  );
  DFFSR _13347_ (
    .CLK(dco_clk),
    .D(_04544_),
    .Q( multiplier_0.reshi_6_ ),
    .R(_04476_),
    .S(1'h1)
  );
  DFFSR _13348_ (
    .CLK(dco_clk),
    .D(_04545_),
    .Q( multiplier_0.reshi_7_ ),
    .R(_04477_),
    .S(1'h1)
  );
  DFFSR _13349_ (
    .CLK(dco_clk),
    .D(_04546_),
    .Q( multiplier_0.reshi_8_ ),
    .R(_04478_),
    .S(1'h1)
  );
  DFFSR _13350_ (
    .CLK(dco_clk),
    .D(_04547_),
    .Q( multiplier_0.reshi_9_ ),
    .R(_04479_),
    .S(1'h1)
  );
  DFFSR _13351_ (
    .CLK(dco_clk),
    .D(_04548_),
    .Q( multiplier_0.reshi_10_ ),
    .R(_04480_),
    .S(1'h1)
  );
  DFFSR _13352_ (
    .CLK(dco_clk),
    .D(_04549_),
    .Q( multiplier_0.reshi_11_ ),
    .R(_04481_),
    .S(1'h1)
  );
  DFFSR _13353_ (
    .CLK(dco_clk),
    .D(_04550_),
    .Q( multiplier_0.reshi_12_ ),
    .R(_04482_),
    .S(1'h1)
  );
  DFFSR _13354_ (
    .CLK(dco_clk),
    .D(_04551_),
    .Q( multiplier_0.reshi_13_ ),
    .R(_04483_),
    .S(1'h1)
  );
  DFFSR _13355_ (
    .CLK(dco_clk),
    .D(_04552_),
    .Q( multiplier_0.reshi_14_ ),
    .R(_04484_),
    .S(1'h1)
  );
  DFFSR _13356_ (
    .CLK(dco_clk),
    .D(_04553_),
    .Q( multiplier_0.reshi_15_ ),
    .R(_04485_),
    .S(1'h1)
  );
  DFFSR _13357_ (
    .CLK(dco_clk),
    .D(_04554_),
    .Q( multiplier_0.reslo_0_ ),
    .R(_04486_),
    .S(1'h1)
  );
  DFFSR _13358_ (
    .CLK(dco_clk),
    .D(_04555_),
    .Q( multiplier_0.reslo_1_ ),
    .R(_04487_),
    .S(1'h1)
  );
  DFFSR _13359_ (
    .CLK(dco_clk),
    .D(_04556_),
    .Q( multiplier_0.reslo_2_ ),
    .R(_04488_),
    .S(1'h1)
  );
  DFFSR _13360_ (
    .CLK(dco_clk),
    .D(_04557_),
    .Q( multiplier_0.reslo_3_ ),
    .R(_04489_),
    .S(1'h1)
  );
  DFFSR _13361_ (
    .CLK(dco_clk),
    .D(_04558_),
    .Q( multiplier_0.reslo_4_ ),
    .R(_04490_),
    .S(1'h1)
  );
  DFFSR _13362_ (
    .CLK(dco_clk),
    .D(_04559_),
    .Q( multiplier_0.reslo_5_ ),
    .R(_04491_),
    .S(1'h1)
  );
  DFFSR _13363_ (
    .CLK(dco_clk),
    .D(_04560_),
    .Q( multiplier_0.reslo_6_ ),
    .R(_04492_),
    .S(1'h1)
  );
  DFFSR _13364_ (
    .CLK(dco_clk),
    .D(_04561_),
    .Q( multiplier_0.reslo_7_ ),
    .R(_04493_),
    .S(1'h1)
  );
  DFFSR _13365_ (
    .CLK(dco_clk),
    .D(_04562_),
    .Q( multiplier_0.reslo_8_ ),
    .R(_04494_),
    .S(1'h1)
  );
  DFFSR _13366_ (
    .CLK(dco_clk),
    .D(_04563_),
    .Q( multiplier_0.reslo_9_ ),
    .R(_04495_),
    .S(1'h1)
  );
  DFFSR _13367_ (
    .CLK(dco_clk),
    .D(_04564_),
    .Q( multiplier_0.reslo_10_ ),
    .R(_04496_),
    .S(1'h1)
  );
  DFFSR _13368_ (
    .CLK(dco_clk),
    .D(_04565_),
    .Q( multiplier_0.reslo_11_ ),
    .R(_04497_),
    .S(1'h1)
  );
  DFFSR _13369_ (
    .CLK(dco_clk),
    .D(_04566_),
    .Q( multiplier_0.reslo_12_ ),
    .R(_04498_),
    .S(1'h1)
  );
  DFFSR _13370_ (
    .CLK(dco_clk),
    .D(_04567_),
    .Q( multiplier_0.reslo_13_ ),
    .R(_04499_),
    .S(1'h1)
  );
  DFFSR _13371_ (
    .CLK(dco_clk),
    .D(_04568_),
    .Q( multiplier_0.reslo_14_ ),
    .R(_04500_),
    .S(1'h1)
  );
  DFFSR _13372_ (
    .CLK(dco_clk),
    .D(_04569_),
    .Q( multiplier_0.reslo_15_ ),
    .R(_04501_),
    .S(1'h1)
  );
  DFFSR _13373_ (
    .CLK(dco_clk),
    .D(_04570_),
    .Q( multiplier_0.op2_0_ ),
    .R(_04502_),
    .S(1'h1)
  );
  DFFSR _13374_ (
    .CLK(dco_clk),
    .D(_04571_),
    .Q( multiplier_0.op2_1_ ),
    .R(_04503_),
    .S(1'h1)
  );
  DFFSR _13375_ (
    .CLK(dco_clk),
    .D(_04572_),
    .Q( multiplier_0.op2_2_ ),
    .R(_04504_),
    .S(1'h1)
  );
  DFFSR _13376_ (
    .CLK(dco_clk),
    .D(_04573_),
    .Q( multiplier_0.op2_3_ ),
    .R(_04505_),
    .S(1'h1)
  );
  DFFSR _13377_ (
    .CLK(dco_clk),
    .D(_04574_),
    .Q( multiplier_0.op2_4_ ),
    .R(_04506_),
    .S(1'h1)
  );
  DFFSR _13378_ (
    .CLK(dco_clk),
    .D(_04575_),
    .Q( multiplier_0.op2_5_ ),
    .R(_04507_),
    .S(1'h1)
  );
  DFFSR _13379_ (
    .CLK(dco_clk),
    .D(_04576_),
    .Q( multiplier_0.op2_6_ ),
    .R(_04508_),
    .S(1'h1)
  );
  DFFSR _13380_ (
    .CLK(dco_clk),
    .D(_04577_),
    .Q( multiplier_0.op2_7_ ),
    .R(_04509_),
    .S(1'h1)
  );
  DFFSR _13381_ (
    .CLK(dco_clk),
    .D(_04578_),
    .Q( multiplier_0.op2_8_ ),
    .R(_04510_),
    .S(1'h1)
  );
  DFFSR _13382_ (
    .CLK(dco_clk),
    .D(_04579_),
    .Q( multiplier_0.op2_9_ ),
    .R(_04511_),
    .S(1'h1)
  );
  DFFSR _13383_ (
    .CLK(dco_clk),
    .D(_04580_),
    .Q( multiplier_0.op2_10_ ),
    .R(_04512_),
    .S(1'h1)
  );
  DFFSR _13384_ (
    .CLK(dco_clk),
    .D(_04581_),
    .Q( multiplier_0.op2_11_ ),
    .R(_04513_),
    .S(1'h1)
  );
  DFFSR _13385_ (
    .CLK(dco_clk),
    .D(_04582_),
    .Q( multiplier_0.op2_12_ ),
    .R(_04514_),
    .S(1'h1)
  );
  DFFSR _13386_ (
    .CLK(dco_clk),
    .D(_04583_),
    .Q( multiplier_0.op2_13_ ),
    .R(_04515_),
    .S(1'h1)
  );
  DFFSR _13387_ (
    .CLK(dco_clk),
    .D(_04584_),
    .Q( multiplier_0.op2_14_ ),
    .R(_04516_),
    .S(1'h1)
  );
  DFFSR _13388_ (
    .CLK(dco_clk),
    .D(_04585_),
    .Q( multiplier_0.op2_15_ ),
    .R(_04517_),
    .S(1'h1)
  );
  DFFSR _13389_ (
    .CLK(dco_clk),
    .D(_04586_),
    .Q( multiplier_0.op1_0_ ),
    .R(_04518_),
    .S(1'h1)
  );
  DFFSR _13390_ (
    .CLK(dco_clk),
    .D(_04587_),
    .Q( multiplier_0.op1_1_ ),
    .R(_04519_),
    .S(1'h1)
  );
  DFFSR _13391_ (
    .CLK(dco_clk),
    .D(_04588_),
    .Q( multiplier_0.op1_2_ ),
    .R(_04520_),
    .S(1'h1)
  );
  DFFSR _13392_ (
    .CLK(dco_clk),
    .D(_04589_),
    .Q( multiplier_0.op1_3_ ),
    .R(_04521_),
    .S(1'h1)
  );
  DFFSR _13393_ (
    .CLK(dco_clk),
    .D(_04590_),
    .Q( multiplier_0.op1_4_ ),
    .R(_04522_),
    .S(1'h1)
  );
  DFFSR _13394_ (
    .CLK(dco_clk),
    .D(_04591_),
    .Q( multiplier_0.op1_5_ ),
    .R(_04523_),
    .S(1'h1)
  );
  DFFSR _13395_ (
    .CLK(dco_clk),
    .D(_04592_),
    .Q( multiplier_0.op1_6_ ),
    .R(_04524_),
    .S(1'h1)
  );
  DFFSR _13396_ (
    .CLK(dco_clk),
    .D(_04593_),
    .Q( multiplier_0.op1_7_ ),
    .R(_04525_),
    .S(1'h1)
  );
  DFFSR _13397_ (
    .CLK(dco_clk),
    .D(_04594_),
    .Q( multiplier_0.op1_8_ ),
    .R(_04526_),
    .S(1'h1)
  );
  DFFSR _13398_ (
    .CLK(dco_clk),
    .D(_04595_),
    .Q( multiplier_0.op1_9_ ),
    .R(_04527_),
    .S(1'h1)
  );
  DFFSR _13399_ (
    .CLK(dco_clk),
    .D(_04596_),
    .Q( multiplier_0.op1_10_ ),
    .R(_04528_),
    .S(1'h1)
  );
  DFFSR _13400_ (
    .CLK(dco_clk),
    .D(_04597_),
    .Q( multiplier_0.op1_11_ ),
    .R(_04529_),
    .S(1'h1)
  );
  DFFSR _13401_ (
    .CLK(dco_clk),
    .D(_04598_),
    .Q( multiplier_0.op1_12_ ),
    .R(_04530_),
    .S(1'h1)
  );
  DFFSR _13402_ (
    .CLK(dco_clk),
    .D(_04599_),
    .Q( multiplier_0.op1_13_ ),
    .R(_04531_),
    .S(1'h1)
  );
  DFFSR _13403_ (
    .CLK(dco_clk),
    .D(_04600_),
    .Q( multiplier_0.op1_14_ ),
    .R(_04532_),
    .S(1'h1)
  );
  DFFSR _13404_ (
    .CLK(dco_clk),
    .D(_04601_),
    .Q( multiplier_0.op1_15_ ),
    .R(_04533_),
    .S(1'h1)
  );
  INVX1 _13405_ (
    .A( sfr_0.ie1_0_ ),
    .Y(_06010_)
  );
  INVX1 _13406_ (
    .A(_06275_),
    .Y(_06011_)
  );
  INVX1 _13407_ (
    .A(_06267_),
    .Y(_06012_)
  );
  INVX1 _13408_ (
    .A(_06265_),
    .Y(_06013_)
  );
  INVX1 _13409_ (
    .A(_06291_),
    .Y(_06014_)
  );
  INVX1 _13410_ (
    .A(1'h0),
    .Y(_06015_)
  );
  INVX1 _13411_ (
    .A(1'h0),
    .Y(_06016_)
  );
  INVX1 _13412_ (
    .A(1'h0),
    .Y(_06017_)
  );
  INVX1 _13413_ (
    .A(1'h0),
    .Y(_06018_)
  );
  INVX1 _13414_ (
    .A(_06327_),
    .Y(_06004_)
  );
  OR2X1 _13415_ (
    .A(_06267_),
    .B(_06262_),
    .Y(_06019_)
  );
  NOR2X1 _13416_ (
    .A(_06266_),
    .B(_06019_),
    .Y(_06020_)
  );
  NOR2X1 _13417_ (
    .A(_06264_),
    .B(1'h0),
    .Y(_06021_)
  );
  OR2X1 _13418_ (
    .A(_06264_),
    .B(1'h0),
    .Y(_06022_)
  );
  NOR3X1 _13419_ (
    .A(_06265_),
    .B(_06014_),
    .C(_06022_),
    .Y(_06023_)
  );
  NAND3X1 _13420_ (
    .A(_06013_),
    .B(_06291_),
    .C(_06021_),
    .Y(_06024_)
  );
  NOR2X1 _13421_ (
    .A(_06273_),
    .B(_06272_),
    .Y(_06025_)
  );
  NOR2X1 _13422_ (
    .A(_06263_),
    .B(_06274_),
    .Y(_06026_)
  );
  AND2X1 _13423_ (
    .A(_06025_),
    .B(_06026_),
    .Y(_06027_)
  );
  NAND2X1 _13424_ (
    .A(_06025_),
    .B(_06026_),
    .Y(_06028_)
  );
  NOR2X1 _13425_ (
    .A(_06269_),
    .B(_06268_),
    .Y(_06029_)
  );
  NOR2X1 _13426_ (
    .A(_06271_),
    .B(_06270_),
    .Y(_06030_)
  );
  AND2X1 _13427_ (
    .A(_06029_),
    .B(_06030_),
    .Y(_06031_)
  );
  NAND2X1 _13428_ (
    .A(_06029_),
    .B(_06030_),
    .Y(_06032_)
  );
  NOR3X1 _13429_ (
    .A(_06024_),
    .B(_06028_),
    .C(_06032_),
    .Y(_06033_)
  );
  NAND3X1 _13430_ (
    .A(_06023_),
    .B(_06027_),
    .C(_06031_),
    .Y(_06034_)
  );
  NAND3X1 _13431_ (
    .A(_06292_),
    .B(_06020_),
    .C(_06033_),
    .Y(_06035_)
  );
  MUX2X1 _13432_ (
    .A(_06010_),
    .B(_06011_),
    .S(_06035_),
    .Y(_06005_)
  );
  NOR2X1 _13433_ (
    .A(_06293_),
    .B(_06292_),
    .Y(_06036_)
  );
  INVX1 _13434_ (
    .A(_06036_),
    .Y(_06037_)
  );
  NAND2X1 _13435_ (
    .A(_06033_),
    .B(_06036_),
    .Y(_06038_)
  );
  NOR3X1 _13436_ (
    .A(_06012_),
    .B(_06262_),
    .C(_06266_),
    .Y(_06039_)
  );
  INVX1 _13437_ (
    .A(_06039_),
    .Y(_06040_)
  );
  NOR3X1 _13438_ (
    .A(_06034_),
    .B(_06037_),
    .C(_06040_),
    .Y(_06041_)
  );
  NAND3X1 _13439_ (
    .A(_06033_),
    .B(_06036_),
    .C(_06039_),
    .Y(_06042_)
  );
  NAND3X1 _13440_ (
    .A(_06266_),
    .B(_06033_),
    .C(_06036_),
    .Y(_06043_)
  );
  OAI22X1 _13441_ (
    .A(_06015_),
    .B(_06042_),
    .C(_06043_),
    .D(_06019_),
    .Y( sfr_0.per_dout_14_ )
  );
  NAND2X1 _13442_ (
    .A(_06012_),
    .B(_06262_),
    .Y(_06044_)
  );
  OAI22X1 _13443_ (
    .A(_06016_),
    .B(_06042_),
    .C(_06043_),
    .D(_06044_),
    .Y( sfr_0.per_dout_8_ )
  );
  OAI22X1 _13444_ (
    .A(_06017_),
    .B(_06042_),
    .C(_06043_),
    .D(_06044_),
    .Y( sfr_0.per_dout_15_ )
  );
  OAI22X1 _13445_ (
    .A(_06018_),
    .B(_06042_),
    .C(_06043_),
    .D(_06019_),
    .Y( sfr_0.per_dout_1_ )
  );
  NOR2X1 _13446_ (
    .A(_06266_),
    .B(_06044_),
    .Y(_06045_)
  );
  NOR2X1 _13447_ (
    .A(_06010_),
    .B(_06262_),
    .Y(_06006_)
  );
  OAI21X1 _13448_ (
    .A(_06266_),
    .B(_06006_),
    .C(_06012_),
    .Y(_06007_)
  );
  AOI22X1 _13449_ (
    .A(1'h0),
    .B(_06039_),
    .C(_06045_),
    .D( sfr_0.ifg1_0_ ),
    .Y(_06008_)
  );
  AOI21X1 _13450_ (
    .A(_06007_),
    .B(_06008_),
    .C(_06038_),
    .Y( sfr_0.per_dout_0_ )
  );
  NAND3X1 _13451_ (
    .A(_06292_),
    .B(_06033_),
    .C(_06045_),
    .Y(_06009_)
  );
  NOR2X1 _13452_ (
    .A(_06275_),
    .B(_06009_),
    .Y( sfr_0.wdtifg_sw_clr )
  );
  NOR2X1 _13453_ (
    .A(_06011_),
    .B(_06009_),
    .Y( sfr_0.wdtifg_sw_set )
  );
  AND2X1 _13454_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_2_ )
  );
  AND2X1 _13455_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_3_ )
  );
  AND2X1 _13456_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_4_ )
  );
  AND2X1 _13457_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_5_ )
  );
  AND2X1 _13458_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_6_ )
  );
  AND2X1 _13459_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_7_ )
  );
  AND2X1 _13460_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_9_ )
  );
  AND2X1 _13461_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_10_ )
  );
  AND2X1 _13462_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_11_ )
  );
  AND2X1 _13463_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_12_ )
  );
  AND2X1 _13464_ (
    .A(1'h0),
    .B(_06041_),
    .Y( sfr_0.cpu_nr_rd_13_ )
  );
  DFFSR _13465_ (
    .CLK(dco_clk),
    .D(_06005_),
    .Q( sfr_0.ie1_0_ ),
    .R(_06004_),
    .S(1'h1)
  );
  INVX1 _13466_ (
    .A( watchdog_0.wdtcnt_13_ ),
    .Y(_06092_)
  );
  INVX1 _13467_ (
    .A( watchdog_0.wdtcnt_11_ ),
    .Y(_06093_)
  );
  INVX1 _13468_ (
    .A( watchdog_0.wdtcnt_10_ ),
    .Y(_06094_)
  );
  INVX1 _13469_ (
    .A( watchdog_0.wdtcnt_9_ ),
    .Y(_06095_)
  );
  INVX1 _13470_ (
    .A( watchdog_0.wdtcnt_8_ ),
    .Y(_06096_)
  );
  INVX1 _13471_ (
    .A( watchdog_0.wdtcnt_7_ ),
    .Y(_06097_)
  );
  INVX1 _13472_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .Y(_06098_)
  );
  INVX1 _13473_ (
    .A( watchdog_0.wdtcnt_2_ ),
    .Y(_06099_)
  );
  INVX1 _13474_ (
    .A( watchdog_0.wdtctl_1_ ),
    .Y(_06100_)
  );
  INVX1 _13475_ (
    .A(_06271_),
    .Y(_06101_)
  );
  INVX1 _13476_ (
    .A(_06273_),
    .Y(_06102_)
  );
  INVX1 _13477_ (
    .A(_06263_),
    .Y(_06103_)
  );
  INVX1 _13478_ (
    .A(_06265_),
    .Y(_06104_)
  );
  INVX1 _13479_ (
    .A(_06291_),
    .Y(_06105_)
  );
  INVX1 _13480_ (
    .A( sfr_0.wdtifg_sw_set ),
    .Y(_06106_)
  );
  INVX1 _13481_ (
    .A( sfr_0.wdtifg_sw_clr ),
    .Y(_06107_)
  );
  INVX1 _13482_ (
    .A( clock_module_0.por ),
    .Y(_06047_)
  );
  INVX1 _13483_ (
    .A(_06327_),
    .Y(_06048_)
  );
  MUX2X1 _13484_ (
    .A(_06213_),
    .B(_06328_),
    .S( watchdog_0.wdtctl_2_ ),
    .Y(_06108_)
  );
  OR2X1 _13485_ (
    .A( watchdog_0.wdtctl_7_ ),
    .B(_06214_),
    .Y(_06109_)
  );
  NOR2X1 _13486_ (
    .A(_06108_),
    .B(_06109_),
    .Y(_06110_)
  );
  INVX1 _13487_ (
    .A(_06110_),
    .Y(_06111_)
  );
  NAND3X1 _13488_ (
    .A( watchdog_0.wdtcnt_5_ ),
    .B( watchdog_0.wdtcnt_2_ ),
    .C( watchdog_0.wdtcnt_0_ ),
    .Y(_06112_)
  );
  NAND3X1 _13489_ (
    .A( watchdog_0.wdtcnt_4_ ),
    .B( watchdog_0.wdtcnt_3_ ),
    .C( watchdog_0.wdtcnt_1_ ),
    .Y(_06113_)
  );
  NOR2X1 _13490_ (
    .A(_06112_),
    .B(_06113_),
    .Y(_06114_)
  );
  NOR3X1 _13491_ (
    .A(_06098_),
    .B(_06112_),
    .C(_06113_),
    .Y(_06115_)
  );
  NOR2X1 _13492_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_06114_),
    .Y(_06116_)
  );
  NOR2X1 _13493_ (
    .A(_06115_),
    .B(_06116_),
    .Y(_06117_)
  );
  NAND3X1 _13494_ (
    .A( watchdog_0.wdtctl_1_ ),
    .B( watchdog_0.wdtctl_0_ ),
    .C(_06117_),
    .Y(_06118_)
  );
  NOR2X1 _13495_ (
    .A( watchdog_0.wdtctl_1_ ),
    .B( watchdog_0.wdtctl_0_ ),
    .Y(_06119_)
  );
  NOR2X1 _13496_ (
    .A(_06096_),
    .B(_06097_),
    .Y(_06120_)
  );
  NAND2X1 _13497_ (
    .A( watchdog_0.wdtcnt_8_ ),
    .B( watchdog_0.wdtcnt_7_ ),
    .Y(_06121_)
  );
  NAND3X1 _13498_ (
    .A( watchdog_0.wdtcnt_9_ ),
    .B(_06115_),
    .C(_06120_),
    .Y(_06122_)
  );
  NAND2X1 _13499_ (
    .A( watchdog_0.wdtcnt_11_ ),
    .B( watchdog_0.wdtcnt_10_ ),
    .Y(_06123_)
  );
  NAND3X1 _13500_ (
    .A( watchdog_0.wdtcnt_12_ ),
    .B( watchdog_0.wdtcnt_11_ ),
    .C( watchdog_0.wdtcnt_10_ ),
    .Y(_06124_)
  );
  NOR2X1 _13501_ (
    .A(_06122_),
    .B(_06124_),
    .Y(_06125_)
  );
  NOR3X1 _13502_ (
    .A(_06092_),
    .B(_06122_),
    .C(_06124_),
    .Y(_06126_)
  );
  NAND2X1 _13503_ (
    .A( watchdog_0.wdtcnt_13_ ),
    .B(_06125_),
    .Y(_06127_)
  );
  OAI21X1 _13504_ (
    .A(_06122_),
    .B(_06124_),
    .C(_06092_),
    .Y(_06128_)
  );
  AND2X1 _13505_ (
    .A(_06100_),
    .B(_06128_),
    .Y(_06129_)
  );
  AOI21X1 _13506_ (
    .A(_06115_),
    .B(_06120_),
    .C( watchdog_0.wdtcnt_9_ ),
    .Y(_06130_)
  );
  NOR2X1 _13507_ (
    .A( watchdog_0.wdtctl_0_ ),
    .B(_06130_),
    .Y(_06131_)
  );
  AOI22X1 _13508_ (
    .A(_06127_),
    .B(_06129_),
    .C(_06131_),
    .D(_06122_),
    .Y(_06132_)
  );
  OAI21X1 _13509_ (
    .A(_06119_),
    .B(_06132_),
    .C(_06118_),
    .Y(_06133_)
  );
  NAND2X1 _13510_ (
    .A(_06110_),
    .B(_06133_),
    .Y(_06134_)
  );
  AND2X1 _13511_ (
    .A( watchdog_0.wdtcnt_14_ ),
    .B(_06126_),
    .Y(_06135_)
  );
  OR2X1 _13512_ (
    .A( watchdog_0.wdtcnt_15_ ),
    .B(_06135_),
    .Y(_06136_)
  );
  AOI21X1 _13513_ (
    .A( watchdog_0.wdtcnt_15_ ),
    .B(_06135_),
    .C(_06111_),
    .Y(_06137_)
  );
  NAND3X1 _13514_ (
    .A(_06119_),
    .B(_06136_),
    .C(_06137_),
    .Y(_06138_)
  );
  OR2X1 _13515_ (
    .A(_06279_),
    .B(_06281_),
    .Y(_06139_)
  );
  NAND2X1 _13516_ (
    .A(_06290_),
    .B(_06277_),
    .Y(_06140_)
  );
  NOR2X1 _13517_ (
    .A(_06289_),
    .B(_06276_),
    .Y(_06141_)
  );
  NAND3X1 _13518_ (
    .A(_06278_),
    .B(_06280_),
    .C(_06141_),
    .Y(_06142_)
  );
  OR2X1 _13519_ (
    .A(_06140_),
    .B(_06142_),
    .Y(_06143_)
  );
  NOR2X1 _13520_ (
    .A(_06293_),
    .B(_06292_),
    .Y(_06144_)
  );
  NOR2X1 _13521_ (
    .A(_06270_),
    .B(_06273_),
    .Y(_06145_)
  );
  NAND3X1 _13522_ (
    .A(_06269_),
    .B(_06101_),
    .C(_06145_),
    .Y(_06146_)
  );
  NOR2X1 _13523_ (
    .A(_06262_),
    .B(_06267_),
    .Y(_06147_)
  );
  NOR2X1 _13524_ (
    .A(_06266_),
    .B(_06268_),
    .Y(_06148_)
  );
  NAND2X1 _13525_ (
    .A(_06147_),
    .B(_06148_),
    .Y(_06149_)
  );
  NOR2X1 _13526_ (
    .A(_06146_),
    .B(_06149_),
    .Y(_06150_)
  );
  NOR2X1 _13527_ (
    .A(_06264_),
    .B(1'h0),
    .Y(_06151_)
  );
  NAND2X1 _13528_ (
    .A(_06291_),
    .B(_06151_),
    .Y(_06152_)
  );
  NOR2X1 _13529_ (
    .A(_06274_),
    .B(_06265_),
    .Y(_06153_)
  );
  NAND3X1 _13530_ (
    .A(_06272_),
    .B(_06103_),
    .C(_06153_),
    .Y(_06154_)
  );
  NOR2X1 _13531_ (
    .A(_06152_),
    .B(_06154_),
    .Y(_06155_)
  );
  NOR2X1 _13532_ (
    .A(_06271_),
    .B(_06270_),
    .Y(_06156_)
  );
  NOR2X1 _13533_ (
    .A(_06262_),
    .B(_06268_),
    .Y(_06157_)
  );
  AND2X1 _13534_ (
    .A(_06156_),
    .B(_06157_),
    .Y(_06158_)
  );
  OR2X1 _13535_ (
    .A(_06263_),
    .B(_06274_),
    .Y(_06159_)
  );
  NOR2X1 _13536_ (
    .A(_06264_),
    .B(_06159_),
    .Y(_06160_)
  );
  NOR2X1 _13537_ (
    .A(_06267_),
    .B(_06266_),
    .Y(_06161_)
  );
  NAND3X1 _13538_ (
    .A(_06269_),
    .B(_06102_),
    .C(_06161_),
    .Y(_06162_)
  );
  NOR2X1 _13539_ (
    .A(1'h0),
    .B(_06105_),
    .Y(_06163_)
  );
  NAND3X1 _13540_ (
    .A(_06272_),
    .B(_06104_),
    .C(_06163_),
    .Y(_06164_)
  );
  NOR2X1 _13541_ (
    .A(_06162_),
    .B(_06164_),
    .Y(_06165_)
  );
  NAND3X1 _13542_ (
    .A(_06158_),
    .B(_06160_),
    .C(_06165_),
    .Y(_06166_)
  );
  NOR2X1 _13543_ (
    .A(_06144_),
    .B(_06166_),
    .Y(_06167_)
  );
  OAI21X1 _13544_ (
    .A(_06139_),
    .B(_06143_),
    .C(_06167_),
    .Y(_06168_)
  );
  AND2X1 _13545_ (
    .A(_06138_),
    .B(_06168_),
    .Y(_06169_)
  );
  AND2X1 _13546_ (
    .A(_06134_),
    .B(_06169_),
    .Y(_06170_)
  );
  NAND2X1 _13547_ (
    .A(_06284_),
    .B(_06167_),
    .Y(_06171_)
  );
  NAND3X1 _13548_ (
    .A(_06134_),
    .B(_06169_),
    .C(_06171_),
    .Y(_06172_)
  );
  AOI22X1 _13549_ (
    .A( watchdog_0.wdtcnt_15_ ),
    .B(_06111_),
    .C(_06136_),
    .D(_06137_),
    .Y(_06173_)
  );
  NOR2X1 _13550_ (
    .A(_06172_),
    .B(_06173_),
    .Y(_06091_)
  );
  NAND2X1 _13551_ (
    .A(_06110_),
    .B(_06125_),
    .Y(_06174_)
  );
  NOR2X1 _13552_ (
    .A(_06111_),
    .B(_06127_),
    .Y(_06175_)
  );
  XNOR2X1 _13553_ (
    .A( watchdog_0.wdtcnt_14_ ),
    .B(_06175_),
    .Y(_06176_)
  );
  NOR2X1 _13554_ (
    .A(_06172_),
    .B(_06176_),
    .Y(_06090_)
  );
  OR2X1 _13555_ (
    .A(_06111_),
    .B(_06122_),
    .Y(_06177_)
  );
  NAND2X1 _13556_ (
    .A(_06110_),
    .B(_06115_),
    .Y(_06178_)
  );
  OAI21X1 _13557_ (
    .A(_06124_),
    .B(_06177_),
    .C(_06092_),
    .Y(_06179_)
  );
  OAI21X1 _13558_ (
    .A(_06111_),
    .B(_06127_),
    .C(_06179_),
    .Y(_06180_)
  );
  NOR2X1 _13559_ (
    .A(_06172_),
    .B(_06180_),
    .Y(_06089_)
  );
  NOR2X1 _13560_ (
    .A(_06123_),
    .B(_06177_),
    .Y(_06181_)
  );
  OAI21X1 _13561_ (
    .A( watchdog_0.wdtcnt_12_ ),
    .B(_06181_),
    .C(_06174_),
    .Y(_06182_)
  );
  NOR2X1 _13562_ (
    .A(_06172_),
    .B(_06182_),
    .Y(_06088_)
  );
  OAI21X1 _13563_ (
    .A(_06094_),
    .B(_06177_),
    .C(_06093_),
    .Y(_06183_)
  );
  OAI21X1 _13564_ (
    .A(_06123_),
    .B(_06177_),
    .C(_06183_),
    .Y(_06184_)
  );
  NOR2X1 _13565_ (
    .A(_06172_),
    .B(_06184_),
    .Y(_06087_)
  );
  XNOR2X1 _13566_ (
    .A(_06094_),
    .B(_06177_),
    .Y(_06185_)
  );
  NOR2X1 _13567_ (
    .A(_06172_),
    .B(_06185_),
    .Y(_06086_)
  );
  OAI21X1 _13568_ (
    .A(_06121_),
    .B(_06178_),
    .C(_06095_),
    .Y(_06186_)
  );
  OAI21X1 _13569_ (
    .A(_06111_),
    .B(_06122_),
    .C(_06186_),
    .Y(_06187_)
  );
  NOR2X1 _13570_ (
    .A(_06172_),
    .B(_06187_),
    .Y(_06085_)
  );
  OAI21X1 _13571_ (
    .A(_06097_),
    .B(_06178_),
    .C(_06096_),
    .Y(_06188_)
  );
  OAI21X1 _13572_ (
    .A(_06121_),
    .B(_06178_),
    .C(_06188_),
    .Y(_06189_)
  );
  NOR2X1 _13573_ (
    .A(_06172_),
    .B(_06189_),
    .Y(_06084_)
  );
  XNOR2X1 _13574_ (
    .A(_06097_),
    .B(_06178_),
    .Y(_06190_)
  );
  NOR2X1 _13575_ (
    .A(_06172_),
    .B(_06190_),
    .Y(_06083_)
  );
  OAI21X1 _13576_ (
    .A(_06108_),
    .B(_06109_),
    .C(_06098_),
    .Y(_06191_)
  );
  OAI21X1 _13577_ (
    .A(_06111_),
    .B(_06117_),
    .C(_06191_),
    .Y(_06192_)
  );
  NOR2X1 _13578_ (
    .A(_06172_),
    .B(_06192_),
    .Y(_06082_)
  );
  NAND2X1 _13579_ (
    .A( watchdog_0.wdtcnt_0_ ),
    .B(_06110_),
    .Y(_06193_)
  );
  NAND3X1 _13580_ (
    .A( watchdog_0.wdtcnt_1_ ),
    .B( watchdog_0.wdtcnt_0_ ),
    .C(_06110_),
    .Y(_06194_)
  );
  NOR2X1 _13581_ (
    .A(_06099_),
    .B(_06194_),
    .Y(_06195_)
  );
  NAND2X1 _13582_ (
    .A( watchdog_0.wdtcnt_3_ ),
    .B(_06195_),
    .Y(_06196_)
  );
  NAND3X1 _13583_ (
    .A( watchdog_0.wdtcnt_4_ ),
    .B( watchdog_0.wdtcnt_3_ ),
    .C(_06195_),
    .Y(_06197_)
  );
  XOR2X1 _13584_ (
    .A( watchdog_0.wdtcnt_5_ ),
    .B(_06197_),
    .Y(_06198_)
  );
  NOR2X1 _13585_ (
    .A(_06172_),
    .B(_06198_),
    .Y(_06081_)
  );
  XOR2X1 _13586_ (
    .A( watchdog_0.wdtcnt_4_ ),
    .B(_06196_),
    .Y(_06199_)
  );
  NOR2X1 _13587_ (
    .A(_06172_),
    .B(_06199_),
    .Y(_06080_)
  );
  XNOR2X1 _13588_ (
    .A( watchdog_0.wdtcnt_3_ ),
    .B(_06195_),
    .Y(_06200_)
  );
  NOR2X1 _13589_ (
    .A(_06172_),
    .B(_06200_),
    .Y(_06079_)
  );
  XNOR2X1 _13590_ (
    .A(_06099_),
    .B(_06194_),
    .Y(_06201_)
  );
  NOR2X1 _13591_ (
    .A(_06172_),
    .B(_06201_),
    .Y(_06078_)
  );
  XOR2X1 _13592_ (
    .A( watchdog_0.wdtcnt_1_ ),
    .B(_06193_),
    .Y(_06202_)
  );
  NOR2X1 _13593_ (
    .A(_06172_),
    .B(_06202_),
    .Y(_06077_)
  );
  XNOR2X1 _13594_ (
    .A( watchdog_0.wdtcnt_0_ ),
    .B(_06110_),
    .Y(_06203_)
  );
  NOR2X1 _13595_ (
    .A(_06172_),
    .B(_06203_),
    .Y(_06076_)
  );
  NAND2X1 _13596_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B(_06249_),
    .Y(_06204_)
  );
  NAND3X1 _13597_ (
    .A( sfr_0.ifg1_0_ ),
    .B(_06107_),
    .C(_06204_),
    .Y(_06205_)
  );
  NAND3X1 _13598_ (
    .A(_06106_),
    .B(_06170_),
    .C(_06205_),
    .Y(_06075_)
  );
  MUX2X1 _13599_ (
    .A(_06288_),
    .B( watchdog_0.wdtctl_7_ ),
    .S(_06167_),
    .Y(_06206_)
  );
  INVX1 _13600_ (
    .A(_06206_),
    .Y(_06074_)
  );
  MUX2X1 _13601_ (
    .A(_06285_),
    .B( watchdog_0.wdtctl_4_ ),
    .S(_06167_),
    .Y(_06207_)
  );
  INVX1 _13602_ (
    .A(_06207_),
    .Y(_06073_)
  );
  MUX2X1 _13603_ (
    .A(_06283_),
    .B( watchdog_0.wdtctl_2_ ),
    .S(_06167_),
    .Y(_06208_)
  );
  INVX1 _13604_ (
    .A(_06208_),
    .Y(_06072_)
  );
  MUX2X1 _13605_ (
    .A(_06282_),
    .B( watchdog_0.wdtctl_1_ ),
    .S(_06167_),
    .Y(_06209_)
  );
  INVX1 _13606_ (
    .A(_06209_),
    .Y(_06071_)
  );
  MUX2X1 _13607_ (
    .A(_06275_),
    .B( watchdog_0.wdtctl_0_ ),
    .S(_06167_),
    .Y(_06210_)
  );
  INVX1 _13608_ (
    .A(_06210_),
    .Y(_06070_)
  );
  NAND3X1 _13609_ (
    .A(_06144_),
    .B(_06150_),
    .C(_06155_),
    .Y(_06211_)
  );
  INVX1 _13610_ (
    .A(_06211_),
    .Y( watchdog_0.per_dout_11_ )
  );
  AND2X1 _13611_ (
    .A( watchdog_0.wdtctl_0_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_0_ )
  );
  NOR2X1 _13612_ (
    .A(_06100_),
    .B(_06211_),
    .Y( watchdog_0.per_dout_1_ )
  );
  AND2X1 _13613_ (
    .A( watchdog_0.wdtctl_2_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_2_ )
  );
  AND2X1 _13614_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_4_ )
  );
  AND2X1 _13615_ (
    .A( watchdog_0.wdtctl_7_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_7_ )
  );
  NAND3X1 _13616_ (
    .A( sfr_0.ifg1_0_ ),
    .B( watchdog_0.wdtctl_4_ ),
    .C( sfr_0.ie1_0_ ),
    .Y(_06212_)
  );
  INVX1 _13617_ (
    .A(_06212_),
    .Y( frontend_0.wdt_irq )
  );
  AOI22X1 _13618_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B(_06168_),
    .C(_06170_),
    .D(_06106_),
    .Y(_06046_)
  );
  INVX1 _13619_ (
    .A(_06327_),
    .Y(_06049_)
  );
  INVX1 _13620_ (
    .A(_06327_),
    .Y(_06050_)
  );
  INVX1 _13621_ (
    .A(_06327_),
    .Y(_06051_)
  );
  INVX1 _13622_ (
    .A(_06327_),
    .Y(_06052_)
  );
  INVX1 _13623_ (
    .A( clock_module_0.por ),
    .Y(_06053_)
  );
  INVX1 _13624_ (
    .A(_06327_),
    .Y(_06054_)
  );
  INVX1 _13625_ (
    .A(_06327_),
    .Y(_06055_)
  );
  INVX1 _13626_ (
    .A(_06327_),
    .Y(_06056_)
  );
  INVX1 _13627_ (
    .A(_06327_),
    .Y(_06057_)
  );
  INVX1 _13628_ (
    .A(_06327_),
    .Y(_06058_)
  );
  INVX1 _13629_ (
    .A(_06327_),
    .Y(_06059_)
  );
  INVX1 _13630_ (
    .A(_06327_),
    .Y(_06060_)
  );
  INVX1 _13631_ (
    .A(_06327_),
    .Y(_06061_)
  );
  INVX1 _13632_ (
    .A(_06327_),
    .Y(_06062_)
  );
  INVX1 _13633_ (
    .A(_06327_),
    .Y(_06063_)
  );
  INVX1 _13634_ (
    .A(_06327_),
    .Y(_06064_)
  );
  INVX1 _13635_ (
    .A(_06327_),
    .Y(_06065_)
  );
  INVX1 _13636_ (
    .A(_06327_),
    .Y(_06066_)
  );
  INVX1 _13637_ (
    .A(_06327_),
    .Y(_06067_)
  );
  INVX1 _13638_ (
    .A(_06327_),
    .Y(_06068_)
  );
  INVX1 _13639_ (
    .A(_06327_),
    .Y(_06069_)
  );
  DFFSR _13640_ (
    .CLK(dco_clk),
    .D(_06046_),
    .Q( clock_module_0.wdt_reset ),
    .R(_06047_),
    .S(1'h1)
  );
  DFFSR _13641_ (
    .CLK(dco_clk),
    .D(_06070_),
    .Q( watchdog_0.wdtctl_0_ ),
    .R(_06048_),
    .S(1'h1)
  );
  DFFSR _13642_ (
    .CLK(dco_clk),
    .D(_06071_),
    .Q( watchdog_0.wdtctl_1_ ),
    .R(_06049_),
    .S(1'h1)
  );
  DFFSR _13643_ (
    .CLK(dco_clk),
    .D(_06072_),
    .Q( watchdog_0.wdtctl_2_ ),
    .R(_06050_),
    .S(1'h1)
  );
  DFFSR _13644_ (
    .CLK(dco_clk),
    .D(_06073_),
    .Q( watchdog_0.wdtctl_4_ ),
    .R(_06051_),
    .S(1'h1)
  );
  DFFSR _13645_ (
    .CLK(dco_clk),
    .D(_06074_),
    .Q( watchdog_0.wdtctl_7_ ),
    .R(_06052_),
    .S(1'h1)
  );
  DFFSR _13646_ (
    .CLK(dco_clk),
    .D(_06075_),
    .Q( sfr_0.ifg1_0_ ),
    .R(_06053_),
    .S(1'h1)
  );
  DFFSR _13647_ (
    .CLK(dco_clk),
    .D(_06076_),
    .Q( watchdog_0.wdtcnt_0_ ),
    .R(_06054_),
    .S(1'h1)
  );
  DFFSR _13648_ (
    .CLK(dco_clk),
    .D(_06077_),
    .Q( watchdog_0.wdtcnt_1_ ),
    .R(_06055_),
    .S(1'h1)
  );
  DFFSR _13649_ (
    .CLK(dco_clk),
    .D(_06078_),
    .Q( watchdog_0.wdtcnt_2_ ),
    .R(_06056_),
    .S(1'h1)
  );
  DFFSR _13650_ (
    .CLK(dco_clk),
    .D(_06079_),
    .Q( watchdog_0.wdtcnt_3_ ),
    .R(_06057_),
    .S(1'h1)
  );
  DFFSR _13651_ (
    .CLK(dco_clk),
    .D(_06080_),
    .Q( watchdog_0.wdtcnt_4_ ),
    .R(_06058_),
    .S(1'h1)
  );
  DFFSR _13652_ (
    .CLK(dco_clk),
    .D(_06081_),
    .Q( watchdog_0.wdtcnt_5_ ),
    .R(_06059_),
    .S(1'h1)
  );
  DFFSR _13653_ (
    .CLK(dco_clk),
    .D(_06082_),
    .Q( watchdog_0.wdtcnt_6_ ),
    .R(_06060_),
    .S(1'h1)
  );
  DFFSR _13654_ (
    .CLK(dco_clk),
    .D(_06083_),
    .Q( watchdog_0.wdtcnt_7_ ),
    .R(_06061_),
    .S(1'h1)
  );
  DFFSR _13655_ (
    .CLK(dco_clk),
    .D(_06084_),
    .Q( watchdog_0.wdtcnt_8_ ),
    .R(_06062_),
    .S(1'h1)
  );
  DFFSR _13656_ (
    .CLK(dco_clk),
    .D(_06085_),
    .Q( watchdog_0.wdtcnt_9_ ),
    .R(_06063_),
    .S(1'h1)
  );
  DFFSR _13657_ (
    .CLK(dco_clk),
    .D(_06086_),
    .Q( watchdog_0.wdtcnt_10_ ),
    .R(_06064_),
    .S(1'h1)
  );
  DFFSR _13658_ (
    .CLK(dco_clk),
    .D(_06087_),
    .Q( watchdog_0.wdtcnt_11_ ),
    .R(_06065_),
    .S(1'h1)
  );
  DFFSR _13659_ (
    .CLK(dco_clk),
    .D(_06088_),
    .Q( watchdog_0.wdtcnt_12_ ),
    .R(_06066_),
    .S(1'h1)
  );
  DFFSR _13660_ (
    .CLK(dco_clk),
    .D(_06089_),
    .Q( watchdog_0.wdtcnt_13_ ),
    .R(_06067_),
    .S(1'h1)
  );
  DFFSR _13661_ (
    .CLK(dco_clk),
    .D(_06090_),
    .Q( watchdog_0.wdtcnt_14_ ),
    .R(_06068_),
    .S(1'h1)
  );
  DFFSR _13662_ (
    .CLK(dco_clk),
    .D(_06091_),
    .Q( watchdog_0.wdtcnt_15_ ),
    .R(_06069_),
    .S(1'h1)
  );
  BUFX2 _13663_ (
    .A(dco_clk),
    .Y(aclk)
  );
  BUFX2 _13664_ (
    .A(_06213_),
    .Y(aclk_en)
  );
  BUFX2 _13665_ (
    .A(_06214_),
    .Y(dbg_freeze)
  );
  BUFX2 _13666_ (
    .A(_06215_),
    .Y(dbg_i2c_sda_out)
  );
  BUFX2 _13667_ (
    .A(1'h1),
    .Y(dbg_uart_txd)
  );
  BUFX2 _13668_ (
    .A(1'h1),
    .Y(dco_enable)
  );
  BUFX2 _13669_ (
    .A(1'h1),
    .Y(dco_wkup)
  );
  BUFX2 _13670_ (
    .A(1'h0),
    .Y(dma_dout_0_)
  );
  BUFX2 _13671_ (
    .A(1'h0),
    .Y(dma_dout_10_)
  );
  BUFX2 _13672_ (
    .A(1'h0),
    .Y(dma_dout_11_)
  );
  BUFX2 _13673_ (
    .A(1'h0),
    .Y(dma_dout_12_)
  );
  BUFX2 _13674_ (
    .A(1'h0),
    .Y(dma_dout_13_)
  );
  BUFX2 _13675_ (
    .A(1'h0),
    .Y(dma_dout_14_)
  );
  BUFX2 _13676_ (
    .A(1'h0),
    .Y(dma_dout_15_)
  );
  BUFX2 _13677_ (
    .A(1'h0),
    .Y(dma_dout_1_)
  );
  BUFX2 _13678_ (
    .A(1'h0),
    .Y(dma_dout_2_)
  );
  BUFX2 _13679_ (
    .A(1'h0),
    .Y(dma_dout_3_)
  );
  BUFX2 _13680_ (
    .A(1'h0),
    .Y(dma_dout_4_)
  );
  BUFX2 _13681_ (
    .A(1'h0),
    .Y(dma_dout_5_)
  );
  BUFX2 _13682_ (
    .A(1'h0),
    .Y(dma_dout_6_)
  );
  BUFX2 _13683_ (
    .A(1'h0),
    .Y(dma_dout_7_)
  );
  BUFX2 _13684_ (
    .A(1'h0),
    .Y(dma_dout_8_)
  );
  BUFX2 _13685_ (
    .A(1'h0),
    .Y(dma_dout_9_)
  );
  BUFX2 _13686_ (
    .A(1'h1),
    .Y(dma_ready)
  );
  BUFX2 _13687_ (
    .A(1'h1),
    .Y(dma_resp)
  );
  BUFX2 _13688_ (
    .A(_06216_),
    .Y(dmem_addr_0_)
  );
  BUFX2 _13689_ (
    .A(_06217_),
    .Y(dmem_addr_10_)
  );
  BUFX2 _13690_ (
    .A(_06218_),
    .Y(dmem_addr_11_)
  );
  BUFX2 _13691_ (
    .A(_06219_),
    .Y(dmem_addr_12_)
  );
  BUFX2 _13692_ (
    .A(_06220_),
    .Y(dmem_addr_1_)
  );
  BUFX2 _13693_ (
    .A(_06221_),
    .Y(dmem_addr_2_)
  );
  BUFX2 _13694_ (
    .A(_06222_),
    .Y(dmem_addr_3_)
  );
  BUFX2 _13695_ (
    .A(_06223_),
    .Y(dmem_addr_4_)
  );
  BUFX2 _13696_ (
    .A(_06224_),
    .Y(dmem_addr_5_)
  );
  BUFX2 _13697_ (
    .A(_06225_),
    .Y(dmem_addr_6_)
  );
  BUFX2 _13698_ (
    .A(_06226_),
    .Y(dmem_addr_7_)
  );
  BUFX2 _13699_ (
    .A(_06227_),
    .Y(dmem_addr_8_)
  );
  BUFX2 _13700_ (
    .A(_06228_),
    .Y(dmem_addr_9_)
  );
  BUFX2 _13701_ (
    .A(_06229_),
    .Y(dmem_cen)
  );
  BUFX2 _13702_ (
    .A(_06230_),
    .Y(dmem_din_0_)
  );
  BUFX2 _13703_ (
    .A(_06231_),
    .Y(dmem_din_10_)
  );
  BUFX2 _13704_ (
    .A(_06232_),
    .Y(dmem_din_11_)
  );
  BUFX2 _13705_ (
    .A(_06233_),
    .Y(dmem_din_12_)
  );
  BUFX2 _13706_ (
    .A(_06234_),
    .Y(dmem_din_13_)
  );
  BUFX2 _13707_ (
    .A(_06235_),
    .Y(dmem_din_14_)
  );
  BUFX2 _13708_ (
    .A(_06236_),
    .Y(dmem_din_15_)
  );
  BUFX2 _13709_ (
    .A(_06237_),
    .Y(dmem_din_1_)
  );
  BUFX2 _13710_ (
    .A(_06238_),
    .Y(dmem_din_2_)
  );
  BUFX2 _13711_ (
    .A(_06239_),
    .Y(dmem_din_3_)
  );
  BUFX2 _13712_ (
    .A(_06240_),
    .Y(dmem_din_4_)
  );
  BUFX2 _13713_ (
    .A(_06241_),
    .Y(dmem_din_5_)
  );
  BUFX2 _13714_ (
    .A(_06242_),
    .Y(dmem_din_6_)
  );
  BUFX2 _13715_ (
    .A(_06243_),
    .Y(dmem_din_7_)
  );
  BUFX2 _13716_ (
    .A(_06244_),
    .Y(dmem_din_8_)
  );
  BUFX2 _13717_ (
    .A(_06245_),
    .Y(dmem_din_9_)
  );
  BUFX2 _13718_ (
    .A(_06246_),
    .Y(dmem_wen_0_)
  );
  BUFX2 _13719_ (
    .A(_06247_),
    .Y(dmem_wen_1_)
  );
  BUFX2 _13720_ (
    .A(_06248_),
    .Y(irq_acc_0_)
  );
  BUFX2 _13721_ (
    .A(_06249_),
    .Y(irq_acc_10_)
  );
  BUFX2 _13722_ (
    .A(_06250_),
    .Y(irq_acc_11_)
  );
  BUFX2 _13723_ (
    .A(_06251_),
    .Y(irq_acc_12_)
  );
  BUFX2 _13724_ (
    .A(_06252_),
    .Y(irq_acc_13_)
  );
  BUFX2 _13725_ (
    .A(_06253_),
    .Y(irq_acc_1_)
  );
  BUFX2 _13726_ (
    .A(_06254_),
    .Y(irq_acc_2_)
  );
  BUFX2 _13727_ (
    .A(_06255_),
    .Y(irq_acc_3_)
  );
  BUFX2 _13728_ (
    .A(_06256_),
    .Y(irq_acc_4_)
  );
  BUFX2 _13729_ (
    .A(_06257_),
    .Y(irq_acc_5_)
  );
  BUFX2 _13730_ (
    .A(_06258_),
    .Y(irq_acc_6_)
  );
  BUFX2 _13731_ (
    .A(_06259_),
    .Y(irq_acc_7_)
  );
  BUFX2 _13732_ (
    .A(_06260_),
    .Y(irq_acc_8_)
  );
  BUFX2 _13733_ (
    .A(_06261_),
    .Y(irq_acc_9_)
  );
  BUFX2 _13734_ (
    .A(1'h1),
    .Y(lfxt_enable)
  );
  BUFX2 _13735_ (
    .A(1'h0),
    .Y(lfxt_wkup)
  );
  BUFX2 _13736_ (
    .A(dco_clk),
    .Y(mclk)
  );
  BUFX2 _13737_ (
    .A(_06262_),
    .Y(per_addr_0_)
  );
  BUFX2 _13738_ (
    .A(_06263_),
    .Y(per_addr_10_)
  );
  BUFX2 _13739_ (
    .A(_06264_),
    .Y(per_addr_11_)
  );
  BUFX2 _13740_ (
    .A(_06265_),
    .Y(per_addr_12_)
  );
  BUFX2 _13741_ (
    .A(1'h0),
    .Y(per_addr_13_)
  );
  BUFX2 _13742_ (
    .A(_06266_),
    .Y(per_addr_1_)
  );
  BUFX2 _13743_ (
    .A(_06267_),
    .Y(per_addr_2_)
  );
  BUFX2 _13744_ (
    .A(_06268_),
    .Y(per_addr_3_)
  );
  BUFX2 _13745_ (
    .A(_06269_),
    .Y(per_addr_4_)
  );
  BUFX2 _13746_ (
    .A(_06270_),
    .Y(per_addr_5_)
  );
  BUFX2 _13747_ (
    .A(_06271_),
    .Y(per_addr_6_)
  );
  BUFX2 _13748_ (
    .A(_06272_),
    .Y(per_addr_7_)
  );
  BUFX2 _13749_ (
    .A(_06273_),
    .Y(per_addr_8_)
  );
  BUFX2 _13750_ (
    .A(_06274_),
    .Y(per_addr_9_)
  );
  BUFX2 _13751_ (
    .A(_06275_),
    .Y(per_din_0_)
  );
  BUFX2 _13752_ (
    .A(_06276_),
    .Y(per_din_10_)
  );
  BUFX2 _13753_ (
    .A(_06277_),
    .Y(per_din_11_)
  );
  BUFX2 _13754_ (
    .A(_06278_),
    .Y(per_din_12_)
  );
  BUFX2 _13755_ (
    .A(_06279_),
    .Y(per_din_13_)
  );
  BUFX2 _13756_ (
    .A(_06280_),
    .Y(per_din_14_)
  );
  BUFX2 _13757_ (
    .A(_06281_),
    .Y(per_din_15_)
  );
  BUFX2 _13758_ (
    .A(_06282_),
    .Y(per_din_1_)
  );
  BUFX2 _13759_ (
    .A(_06283_),
    .Y(per_din_2_)
  );
  BUFX2 _13760_ (
    .A(_06284_),
    .Y(per_din_3_)
  );
  BUFX2 _13761_ (
    .A(_06285_),
    .Y(per_din_4_)
  );
  BUFX2 _13762_ (
    .A(_06286_),
    .Y(per_din_5_)
  );
  BUFX2 _13763_ (
    .A(_06287_),
    .Y(per_din_6_)
  );
  BUFX2 _13764_ (
    .A(_06288_),
    .Y(per_din_7_)
  );
  BUFX2 _13765_ (
    .A(_06289_),
    .Y(per_din_8_)
  );
  BUFX2 _13766_ (
    .A(_06290_),
    .Y(per_din_9_)
  );
  BUFX2 _13767_ (
    .A(_06291_),
    .Y(per_en)
  );
  BUFX2 _13768_ (
    .A(_06292_),
    .Y(per_we_0_)
  );
  BUFX2 _13769_ (
    .A(_06293_),
    .Y(per_we_1_)
  );
  BUFX2 _13770_ (
    .A(_06294_),
    .Y(pmem_addr_0_)
  );
  BUFX2 _13771_ (
    .A(_06295_),
    .Y(pmem_addr_10_)
  );
  BUFX2 _13772_ (
    .A(_06296_),
    .Y(pmem_addr_11_)
  );
  BUFX2 _13773_ (
    .A(_06297_),
    .Y(pmem_addr_12_)
  );
  BUFX2 _13774_ (
    .A(_06298_),
    .Y(pmem_addr_13_)
  );
  BUFX2 _13775_ (
    .A(_06299_),
    .Y(pmem_addr_1_)
  );
  BUFX2 _13776_ (
    .A(_06300_),
    .Y(pmem_addr_2_)
  );
  BUFX2 _13777_ (
    .A(_06301_),
    .Y(pmem_addr_3_)
  );
  BUFX2 _13778_ (
    .A(_06302_),
    .Y(pmem_addr_4_)
  );
  BUFX2 _13779_ (
    .A(_06303_),
    .Y(pmem_addr_5_)
  );
  BUFX2 _13780_ (
    .A(_06304_),
    .Y(pmem_addr_6_)
  );
  BUFX2 _13781_ (
    .A(_06305_),
    .Y(pmem_addr_7_)
  );
  BUFX2 _13782_ (
    .A(_06306_),
    .Y(pmem_addr_8_)
  );
  BUFX2 _13783_ (
    .A(_06307_),
    .Y(pmem_addr_9_)
  );
  BUFX2 _13784_ (
    .A(_06308_),
    .Y(pmem_cen)
  );
  BUFX2 _13785_ (
    .A(_06309_),
    .Y(pmem_din_0_)
  );
  BUFX2 _13786_ (
    .A(_06310_),
    .Y(pmem_din_10_)
  );
  BUFX2 _13787_ (
    .A(_06311_),
    .Y(pmem_din_11_)
  );
  BUFX2 _13788_ (
    .A(_06312_),
    .Y(pmem_din_12_)
  );
  BUFX2 _13789_ (
    .A(_06313_),
    .Y(pmem_din_13_)
  );
  BUFX2 _13790_ (
    .A(_06314_),
    .Y(pmem_din_14_)
  );
  BUFX2 _13791_ (
    .A(_06315_),
    .Y(pmem_din_15_)
  );
  BUFX2 _13792_ (
    .A(_06316_),
    .Y(pmem_din_1_)
  );
  BUFX2 _13793_ (
    .A(_06317_),
    .Y(pmem_din_2_)
  );
  BUFX2 _13794_ (
    .A(_06318_),
    .Y(pmem_din_3_)
  );
  BUFX2 _13795_ (
    .A(_06319_),
    .Y(pmem_din_4_)
  );
  BUFX2 _13796_ (
    .A(_06320_),
    .Y(pmem_din_5_)
  );
  BUFX2 _13797_ (
    .A(_06321_),
    .Y(pmem_din_6_)
  );
  BUFX2 _13798_ (
    .A(_06322_),
    .Y(pmem_din_7_)
  );
  BUFX2 _13799_ (
    .A(_06323_),
    .Y(pmem_din_8_)
  );
  BUFX2 _13800_ (
    .A(_06324_),
    .Y(pmem_din_9_)
  );
  BUFX2 _13801_ (
    .A(_06325_),
    .Y(pmem_wen_0_)
  );
  BUFX2 _13802_ (
    .A(_06326_),
    .Y(pmem_wen_1_)
  );
  BUFX2 _13803_ (
    .A(_06327_),
    .Y(puc_rst)
  );
  BUFX2 _13804_ (
    .A(dco_clk),
    .Y(smclk)
  );
  BUFX2 _13805_ (
    .A(_06328_),
    .Y(smclk_en)
  );
endmodule
